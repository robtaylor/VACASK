.title Top block test simulation
.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.subckt DP8TClockGenerator_8S1R vss vdd clk decodeclk columnclk precharge_n wl_en we_en
Xnonovl vss vdd clk firststage[0] firststage[1] firststage[2] firststage[3] firststage[4] firststage[5] firststage[6] firstpulse firststage[8] secondstage[0] secondstage[1] secondstage[2] secondstage[3] secondstage[4] secondstage[5] secondstage[6] secondpulse secondstage[8] DP8TNonOverlapClock_8S1R
Xdecodeclkbuf vdd vss clk decodeclk buf_x1
Xprechargeinv vdd vss secondpulse precharge_n inv_x1
Xwlenbuf vdd vss firstpulse wl_en buf_x1
Xcolumnclkbuf vdd vss clk columnclk buf_x1
Xweenbuf vdd vss firstpulse we_en buf_x1
.ends DP8TClockGenerator_8S1R

.subckt DP8TLatchedDecoder_2A2R vss vdd clk a[0] a[1] line[0] line[1] line[2] line[3]
Xaff[0] vdd vss a[0] clk aint[0] DP8TDec_dff_x1
Xaff[1] vdd vss a[1] clk aint[1] DP8TDec_dff_x1
Xainv[0] vdd vss aint[0] aint_n[0] DP8TDec_inv_x1
Xainv[1] vdd vss aint[1] aint_n[1] DP8TDec_inv_x1
Xlinenand[0] vdd vss line_n[0] aint_n[0] aint_n[1] DP8TDec_nand2_x0
Xlinenand[1] vdd vss line_n[1] aint[0] aint_n[1] DP8TDec_nand2_x0
Xlinenand[2] vdd vss line_n[2] aint_n[0] aint[1] DP8TDec_nand2_x0
Xlinenand[3] vdd vss line_n[3] aint[0] aint[1] DP8TDec_nand2_x0
Xlineinv[0] vdd vss line_n[0] line[0] DP8TDec_inv_x2
Xlineinv[1] vdd vss line_n[1] line[1] DP8TDec_inv_x2
Xlineinv[2] vdd vss line_n[2] line[2] DP8TDec_inv_x2
Xlineinv[3] vdd vss line_n[3] line[3] DP8TDec_inv_x2
.ends DP8TLatchedDecoder_2A2R

.subckt DP8TDec_dff_x1 vdd vss i clk q
Xclk_nmos _clk_n clk vss vss sg13_lv_nmos l=0.13um w=0.78um
Xclk_pmos _clk_n clk vdd vdd sg13_lv_pmos l=0.13um w=1.2um
Xclk_n_nmos0 vss _clk_n _clk_buf vss sg13_lv_nmos l=0.13um w=0.78um
Xclk_n_pmos0 vdd _clk_n _clk_buf vdd sg13_lv_pmos l=0.13um w=1.2um
Xi_nmos _u i vss vss sg13_lv_nmos l=0.13um w=0.78um
Xi_pmos _u i vdd vdd sg13_lv_pmos l=0.13um w=1.2um
Xu_nmos vss _u _net0 vss sg13_lv_nmos l=0.13um w=0.78um
Xu_pmos vdd _u _net1 vdd sg13_lv_pmos l=0.13um w=1.2um
Xclk_n_nmos1 _net0 _clk_n _dff_m vss sg13_lv_nmos l=0.13um w=0.78um
Xclk_buf_pmos0 _net1 _clk_buf _dff_m vdd sg13_lv_pmos l=0.13um w=1.2um
Xclk_buf_nmos0 _dff_m _clk_buf _net2 vss sg13_lv_nmos l=0.13um w=0.78um
Xclk_n_pmos1 _dff_m _clk_n _net3 vdd sg13_lv_pmos l=0.13um w=1.2um
Xy_nmos _net2 _y vss vss sg13_lv_nmos l=0.13um w=0.78um
Xy_pmos _net3 _y vdd vdd sg13_lv_pmos l=0.13um w=1.2um
Xdff_m_nmos vss _dff_m _y vss sg13_lv_nmos l=0.13um w=0.78um
Xdff_m_pmos vdd _dff_m _y vdd sg13_lv_pmos l=0.13um w=1.2um
Xclk_buf_nmos1 _y _clk_buf _dff_s vss sg13_lv_nmos l=0.13um w=0.78um
Xclk_n_pmos2 _y _clk_n _dff_s vdd sg13_lv_pmos l=0.13um w=1.2um
Xclk_n_nmos2 _dff_s _clk_n _net4 vss sg13_lv_nmos l=0.13um w=0.78um
Xclk_buf_pmos1 _dff_s _clk_buf _net5 vdd sg13_lv_pmos l=0.13um w=1.2um
Xq_nmos _net4 q vss vss sg13_lv_nmos l=0.13um w=0.78um
Xq_pmos _net5 q vdd vdd sg13_lv_pmos l=0.13um w=1.2um
Xdff_s_nmos vss _dff_s q vss sg13_lv_nmos l=0.13um w=2.17um
Xdff_s_pmos vdd _dff_s q vdd sg13_lv_pmos l=0.13um w=3.77um
.ends DP8TDec_dff_x1

.subckt DP8TDec_inv_x1 vdd vss i nq
Xnmos vss i nq vss sg13_lv_nmos l=0.13um w=2.8um
Xpmos vdd i nq vdd sg13_lv_pmos l=0.13um w=4.4um
.ends DP8TDec_inv_x1

.subckt DP8TDec_and3_x1 vdd vss q i0 i1 i2
Xi0_nmos nq i0 _net0 vss sg13_lv_nmos l=0.13um w=0.78um
Xi0_pmos nq i0 vdd vdd sg13_lv_pmos l=0.13um w=1.2um
Xi1_nmos _net0 i1 _net1 vss sg13_lv_nmos l=0.13um w=0.78um
Xi1_pmos vdd i1 nq vdd sg13_lv_pmos l=0.13um w=1.2um
Xi2_nmos _net1 i2 vss vss sg13_lv_nmos l=0.13um w=0.78um
Xi2_pmos nq i2 vdd vdd sg13_lv_pmos l=0.13um w=1.2um
Xn_pd vss nq q vss sg13_lv_nmos l=0.13um w=2.8um
Xq_pu vdd nq q vdd sg13_lv_pmos l=0.13um w=4.4um
.ends DP8TDec_and3_x1

.subckt DP8TDec_and4_x1 vdd vss q i0 i1 i2 i3
Xi0_nmos nq i0 _net0 vss sg13_lv_nmos l=0.13um w=0.78um
Xi0_pmos vdd i0 nq vdd sg13_lv_pmos l=0.13um w=1.2um
Xi1_nmos _net0 i1 _net1 vss sg13_lv_nmos l=0.13um w=0.78um
Xi1_pmos nq i1 vdd vdd sg13_lv_pmos l=0.13um w=1.2um
Xi2_nmos _net1 i2 _net2 vss sg13_lv_nmos l=0.13um w=0.78um
Xi2_pmos vdd i2 nq vdd sg13_lv_pmos l=0.13um w=1.2um
Xi3_nmos _net2 i3 vss vss sg13_lv_nmos l=0.13um w=0.78um
Xi3_pmos nq i3 vdd vdd sg13_lv_pmos l=0.13um w=1.2um
Xn_pd vss nq q vss sg13_lv_nmos l=0.13um w=2.8um
Xq_pu vdd nq q vdd sg13_lv_pmos l=0.13um w=4.4um
.ends DP8TDec_and4_x1

.subckt DP8TRowPredecoders_3_4B_wl1 vss vdd clk a[0] a[1] a[2] a[3] a[4] a[5] a[6] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[0] page[1] page[2] page[3] page[4] page[5] page[6] page[7] page[8] page[9] page[10] page[11] page[12] page[13] page[14] page[15]
Xaff[0] vdd vss a[0] clk aint[0] DP8TDec_dff_x1
Xaff[1] vdd vss a[1] clk aint[1] DP8TDec_dff_x1
Xaff[2] vdd vss a[2] clk aint[2] DP8TDec_dff_x1
Xaff[3] vdd vss a[3] clk aint[3] DP8TDec_dff_x1
Xaff[4] vdd vss a[4] clk aint[4] DP8TDec_dff_x1
Xaff[5] vdd vss a[5] clk aint[5] DP8TDec_dff_x1
Xaff[6] vdd vss a[6] clk aint[6] DP8TDec_dff_x1
Xainv[0] vdd vss aint[0] aint_n[0] DP8TDec_inv_x1
Xainv[1] vdd vss aint[1] aint_n[1] DP8TDec_inv_x1
Xainv[2] vdd vss aint[2] aint_n[2] DP8TDec_inv_x1
Xainv[3] vdd vss aint[3] aint_n[3] DP8TDec_inv_x1
Xainv[4] vdd vss aint[4] aint_n[4] DP8TDec_inv_x1
Xainv[5] vdd vss aint[5] aint_n[5] DP8TDec_inv_x1
Xainv[6] vdd vss aint[6] aint_n[6] DP8TDec_inv_x1
Xpd[0]and[0] vdd vss pd[0][0] aint_n[0] aint_n[1] aint_n[2] DP8TDec_and3_x1
Xpd[0]and[1] vdd vss pd[0][1] aint[0] aint_n[1] aint_n[2] DP8TDec_and3_x1
Xpd[0]and[2] vdd vss pd[0][2] aint_n[0] aint[1] aint_n[2] DP8TDec_and3_x1
Xpd[0]and[3] vdd vss pd[0][3] aint[0] aint[1] aint_n[2] DP8TDec_and3_x1
Xpd[0]and[4] vdd vss pd[0][4] aint_n[0] aint_n[1] aint[2] DP8TDec_and3_x1
Xpd[0]and[5] vdd vss pd[0][5] aint[0] aint_n[1] aint[2] DP8TDec_and3_x1
Xpd[0]and[6] vdd vss pd[0][6] aint_n[0] aint[1] aint[2] DP8TDec_and3_x1
Xpd[0]and[7] vdd vss pd[0][7] aint[0] aint[1] aint[2] DP8TDec_and3_x1
Xpage_and[0] vdd vss page[0] aint_n[3] aint_n[4] aint_n[5] aint_n[6] DP8TDec_and4_x1
Xpage_and[1] vdd vss page[1] aint[3] aint_n[4] aint_n[5] aint_n[6] DP8TDec_and4_x1
Xpage_and[2] vdd vss page[2] aint_n[3] aint[4] aint_n[5] aint_n[6] DP8TDec_and4_x1
Xpage_and[3] vdd vss page[3] aint[3] aint[4] aint_n[5] aint_n[6] DP8TDec_and4_x1
Xpage_and[4] vdd vss page[4] aint_n[3] aint_n[4] aint[5] aint_n[6] DP8TDec_and4_x1
Xpage_and[5] vdd vss page[5] aint[3] aint_n[4] aint[5] aint_n[6] DP8TDec_and4_x1
Xpage_and[6] vdd vss page[6] aint_n[3] aint[4] aint[5] aint_n[6] DP8TDec_and4_x1
Xpage_and[7] vdd vss page[7] aint[3] aint[4] aint[5] aint_n[6] DP8TDec_and4_x1
Xpage_and[8] vdd vss page[8] aint_n[3] aint_n[4] aint_n[5] aint[6] DP8TDec_and4_x1
Xpage_and[9] vdd vss page[9] aint[3] aint_n[4] aint_n[5] aint[6] DP8TDec_and4_x1
Xpage_and[10] vdd vss page[10] aint_n[3] aint[4] aint_n[5] aint[6] DP8TDec_and4_x1
Xpage_and[11] vdd vss page[11] aint[3] aint[4] aint_n[5] aint[6] DP8TDec_and4_x1
Xpage_and[12] vdd vss page[12] aint_n[3] aint_n[4] aint[5] aint[6] DP8TDec_and4_x1
Xpage_and[13] vdd vss page[13] aint[3] aint_n[4] aint[5] aint[6] DP8TDec_and4_x1
Xpage_and[14] vdd vss page[14] aint_n[3] aint[4] aint[5] aint[6] DP8TDec_and4_x1
Xpage_and[15] vdd vss page[15] aint[3] aint[4] aint[5] aint[6] DP8TDec_and4_x1
.ends DP8TRowPredecoders_3_4B_wl1

.subckt DP8TRowDecoderNand3X2 vss vdd pd[0][0] pd[0][1] page wl_en wl_n[0] wl_n[1]
Xnmos[0] wl_n[0] wl_en int[0] vss sg13_lv_nmos l=0.13um w=0.5um
Xnmos[1] int[0] pd[0][0] int[1] vss sg13_lv_nmos l=0.13um w=0.5um
Xnmos[2] int[1] page vss vss sg13_lv_nmos l=0.13um w=0.5um
Xnmos[3] vss page int[2] vss sg13_lv_nmos l=0.13um w=0.5um
Xnmos[4] int[2] pd[0][1] int[3] vss sg13_lv_nmos l=0.13um w=0.5um
Xnmos[5] int[3] wl_en wl_n[1] vss sg13_lv_nmos l=0.13um w=0.5um
Xpmos[0] wl_n[0] wl_en vdd vdd sg13_lv_pmos l=0.13um w=0.5um
Xpmos[1] vdd pd[0][0] wl_n[0] vdd sg13_lv_pmos l=0.13um w=0.5um
Xpmos[2] wl_n[0] page vdd vdd sg13_lv_pmos l=0.13um w=0.5um
Xpmos[3] vdd page wl_n[1] vdd sg13_lv_pmos l=0.13um w=0.5um
Xpmos[4] wl_n[1] pd[0][1] vdd vdd sg13_lv_pmos l=0.13um w=0.5um
Xpmos[5] vdd wl_en wl_n[1] vdd sg13_lv_pmos l=0.13um w=0.5um
.ends DP8TRowDecoderNand3X2

.subckt DP8TWLDrive_26LN100WN26LP200WP_wl1 vss substrate vdd nwell wl_n wl_drive
Xnmos1 vss wl_n wl_drive substrate sg13_lv_nmos l=0.13um w=0.5um
Xnmos2 wl_drive wl_n vss substrate sg13_lv_nmos l=0.13um w=0.5um
Xpmos1 vdd wl_n wl_drive nwell sg13_lv_pmos l=0.13um w=1.0um
Xpmos2 wl_drive wl_n vdd nwell sg13_lv_pmos l=0.13um w=1.0um
.ends DP8TWLDrive_26LN100WN26LP200WP_wl1

.subckt DP8TRowDecoderDriverPage_2PD8R_wl1 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page wl_en
Xnand3[0] vss vdd pd[0][0] pd[0][1] page wl_en wl_n[0] wl_n[1] DP8TRowDecoderNand3X2
Xnand3[1] vss vdd pd[0][2] pd[0][3] page wl_en wl_n[2] wl_n[3] DP8TRowDecoderNand3X2
Xnand3[2] vss vdd pd[0][4] pd[0][5] page wl_en wl_n[4] wl_n[5] DP8TRowDecoderNand3X2
Xnand3[3] vss vdd pd[0][6] pd[0][7] page wl_en wl_n[6] wl_n[7] DP8TRowDecoderNand3X2
Xdrive[0] vss vss vdd vdd wl_n[0] wl[0] DP8TWLDrive_26LN100WN26LP200WP_wl1
Xdrive[1] vss vss vdd vdd wl_n[1] wl[1] DP8TWLDrive_26LN100WN26LP200WP_wl1
Xdrive[2] vss vss vdd vdd wl_n[2] wl[2] DP8TWLDrive_26LN100WN26LP200WP_wl1
Xdrive[3] vss vss vdd vdd wl_n[3] wl[3] DP8TWLDrive_26LN100WN26LP200WP_wl1
Xdrive[4] vss vss vdd vdd wl_n[4] wl[4] DP8TWLDrive_26LN100WN26LP200WP_wl1
Xdrive[5] vss vss vdd vdd wl_n[5] wl[5] DP8TWLDrive_26LN100WN26LP200WP_wl1
Xdrive[6] vss vss vdd vdd wl_n[6] wl[6] DP8TWLDrive_26LN100WN26LP200WP_wl1
Xdrive[7] vss vss vdd vdd wl_n[7] wl[7] DP8TWLDrive_26LN100WN26LP200WP_wl1
.ends DP8TRowDecoderDriverPage_2PD8R_wl1

.subckt DP8TRowDecoderBulkConn vdd vss

.ends DP8TRowDecoderBulkConn

.subckt DP8TRowDecoder_3_4B_wl1 vss vdd a[0] a[1] a[2] a[3] a[4] a[5] a[6] clk wl_en wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127]
Xpredec vss vdd clk a[0] a[1] a[2] a[3] a[4] a[5] a[6] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[0] page[1] page[2] page[3] page[4] page[5] page[6] page[7] page[8] page[9] page[10] page[11] page[12] page[13] page[14] page[15] DP8TRowPredecoders_3_4B_wl1
Xpage[0] vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[0] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[1] vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[1] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[2] vss vdd wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[2] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[3] vss vdd wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[3] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[4] vss vdd wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[4] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[5] vss vdd wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[5] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[6] vss vdd wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[6] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[7] vss vdd wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[7] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[8] vss vdd wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[8] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[9] vss vdd wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[9] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[10] vss vdd wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[10] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[11] vss vdd wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[11] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[12] vss vdd wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[12] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[13] vss vdd wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[13] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[14] vss vdd wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[14] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xpage[15] vss vdd wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[15] wl_en DP8TRowDecoderDriverPage_2PD8R_wl1
Xbulkcon[0] vdd vss DP8TRowDecoderBulkConn
Xbulkcon[1] vdd vss DP8TRowDecoderBulkConn
Xbulkcon[2] vdd vss DP8TRowDecoderBulkConn
Xbulkcon[3] vdd vss DP8TRowDecoderBulkConn
Xbulkcon[4] vdd vss DP8TRowDecoderBulkConn
Xbulkcon[5] vdd vss DP8TRowDecoderBulkConn
Xbulkcon[6] vdd vss DP8TRowDecoderBulkConn
Xbulkcon[7] vdd vss DP8TRowDecoderBulkConn
Xbulkcon[8] vdd vss DP8TRowDecoderBulkConn
.ends DP8TRowDecoder_3_4B_wl1

.subckt DP8TRowPeriphery_3_4_2_wl1 vss vdd clk a[0] a[1] a[2] a[3] a[4] a[5] a[6] a[7] a[8] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] mux[0] mux[1] mux[2] mux[3] columnclk precharge_n we_en
Xclkgen vss vdd clk decodeclk columnclk precharge_n wl_en we_en DP8TClockGenerator_8S1R
Xcoldec vss vdd decodeclk a[0] a[1] mux[0] mux[1] mux[2] mux[3] DP8TLatchedDecoder_2A2R
Xrowdec vss vdd a[2] a[3] a[4] a[5] a[6] a[7] a[8] decodeclk wl_en wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] DP8TRowDecoder_3_4B_wl1
.ends DP8TRowPeriphery_3_4_2_wl1

.subckt nand2_x0 vdd vss nq i0 i1
Xi0_nmos vss i0 _net0 vss sg13_lv_nmos l=0.13um w=0.78um
Xi0_pmos vdd i0 nq vdd sg13_lv_pmos l=0.13um w=0.78um
Xi1_nmos _net0 i1 nq vss sg13_lv_nmos l=0.13um w=0.78um
Xi1_pmos nq i1 vdd vdd sg13_lv_pmos l=0.13um w=0.78um
.ends nand2_x0

.subckt inv_x0 vdd vss i nq
Xnmos vss i nq vss sg13_lv_nmos l=0.13um w=0.78um
Xpmos vdd i nq vdd sg13_lv_pmos l=0.13um w=0.78um
.ends inv_x0

.subckt DP8TNonOverlapClock_8S1R vss vdd clk firststage[0] firststage[1] firststage[2] firststage[3] firststage[4] firststage[5] firststage[6] firststage[7] firststage[8] secondstage[0] secondstage[1] secondstage[2] secondstage[3] secondstage[4] secondstage[5] secondstage[6] secondstage[7] secondstage[8]
Xclkinv vdd vss clk clk_n inv_x0
Xfirstnand2 vdd vss firststage[0] clk secondstage[8] nand2_x0
Xfirststage[0] vdd vss firststage[0] firststage[1] inv_x0
Xfirststage[1] vdd vss firststage[1] firststage[2] inv_x0
Xfirststage[2] vdd vss firststage[2] firststage[3] inv_x0
Xfirststage[3] vdd vss firststage[3] firststage[4] inv_x0
Xfirststage[4] vdd vss firststage[4] firststage[5] inv_x0
Xfirststage[5] vdd vss firststage[5] firststage[6] inv_x0
Xfirststage[6] vdd vss firststage[6] firststage[7] inv_x0
Xfirststage[7] vdd vss firststage[7] firststage[8] inv_x0
Xsecondnand2 vdd vss secondstage[0] clk_n firststage[8] nand2_x0
Xsecondstage[0] vdd vss secondstage[0] secondstage[1] inv_x0
Xsecondstage[1] vdd vss secondstage[1] secondstage[2] inv_x0
Xsecondstage[2] vdd vss secondstage[2] secondstage[3] inv_x0
Xsecondstage[3] vdd vss secondstage[3] secondstage[4] inv_x0
Xsecondstage[4] vdd vss secondstage[4] secondstage[5] inv_x0
Xsecondstage[5] vdd vss secondstage[5] secondstage[6] inv_x0
Xsecondstage[6] vdd vss secondstage[6] secondstage[7] inv_x0
Xsecondstage[7] vdd vss secondstage[7] secondstage[8] inv_x0
.ends DP8TNonOverlapClock_8S1R

.subckt inv_x1 vdd vss i nq
Xnmos vss i nq vss sg13_lv_nmos l=0.13um w=1.46um
Xpmos vdd i nq vdd sg13_lv_pmos l=0.13um w=1.45um
.ends inv_x1

.subckt buf_x1 vdd vss i q
Xstage0_nmos _i_n i vss vss sg13_lv_nmos l=0.13um w=0.78um
Xstage0_pmos _i_n i vdd vdd sg13_lv_pmos l=0.13um w=0.78um
Xnmos vss _i_n q vss sg13_lv_nmos l=0.13um w=1.07um
Xpmos vdd _i_n q vdd sg13_lv_pmos l=0.13um w=1.06um
.ends buf_x1

.subckt DP8TDec_nand2_x0 vdd vss nq i0 i1
Xi0_nmos vss i0 _net0 vss sg13_lv_nmos l=0.13um w=0.78um
Xi0_pmos vdd i0 nq vdd sg13_lv_pmos l=0.13um w=1.2um
Xi1_nmos _net0 i1 nq vss sg13_lv_nmos l=0.13um w=0.78um
Xi1_pmos nq i1 vdd vdd sg13_lv_pmos l=0.13um w=1.2um
.ends DP8TDec_nand2_x0

.subckt DP8TDec_inv_x2 vdd vss i nq
Xnmos[0] vss i nq vss sg13_lv_nmos l=0.13um w=2.8um
Xpmos[0] vdd i nq vdd sg13_lv_pmos l=0.13um w=4.4um
Xnmos[1] nq i vss vss sg13_lv_nmos l=0.13um w=2.8um
Xpmos[1] nq i vdd vdd sg13_lv_pmos l=0.13um w=4.4um
.ends DP8TDec_inv_x2

.subckt DP8TRowPredecoders_3_4B_wl2 vss vdd clk a[0] a[1] a[2] a[3] a[4] a[5] a[6] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[0] page[1] page[2] page[3] page[4] page[5] page[6] page[7] page[8] page[9] page[10] page[11] page[12] page[13] page[14] page[15]
Xaff[0] vdd vss a[0] clk aint[0] DP8TDec_dff_x1
Xaff[1] vdd vss a[1] clk aint[1] DP8TDec_dff_x1
Xaff[2] vdd vss a[2] clk aint[2] DP8TDec_dff_x1
Xaff[3] vdd vss a[3] clk aint[3] DP8TDec_dff_x1
Xaff[4] vdd vss a[4] clk aint[4] DP8TDec_dff_x1
Xaff[5] vdd vss a[5] clk aint[5] DP8TDec_dff_x1
Xaff[6] vdd vss a[6] clk aint[6] DP8TDec_dff_x1
Xainv[0] vdd vss aint[0] aint_n[0] DP8TDec_inv_x1
Xainv[1] vdd vss aint[1] aint_n[1] DP8TDec_inv_x1
Xainv[2] vdd vss aint[2] aint_n[2] DP8TDec_inv_x1
Xainv[3] vdd vss aint[3] aint_n[3] DP8TDec_inv_x1
Xainv[4] vdd vss aint[4] aint_n[4] DP8TDec_inv_x1
Xainv[5] vdd vss aint[5] aint_n[5] DP8TDec_inv_x1
Xainv[6] vdd vss aint[6] aint_n[6] DP8TDec_inv_x1
Xpd[0]and[0] vdd vss pd[0][0] aint_n[0] aint_n[1] aint_n[2] DP8TDec_and3_x1
Xpd[0]and[1] vdd vss pd[0][1] aint[0] aint_n[1] aint_n[2] DP8TDec_and3_x1
Xpd[0]and[2] vdd vss pd[0][2] aint_n[0] aint[1] aint_n[2] DP8TDec_and3_x1
Xpd[0]and[3] vdd vss pd[0][3] aint[0] aint[1] aint_n[2] DP8TDec_and3_x1
Xpd[0]and[4] vdd vss pd[0][4] aint_n[0] aint_n[1] aint[2] DP8TDec_and3_x1
Xpd[0]and[5] vdd vss pd[0][5] aint[0] aint_n[1] aint[2] DP8TDec_and3_x1
Xpd[0]and[6] vdd vss pd[0][6] aint_n[0] aint[1] aint[2] DP8TDec_and3_x1
Xpd[0]and[7] vdd vss pd[0][7] aint[0] aint[1] aint[2] DP8TDec_and3_x1
Xpage_and[0] vdd vss page[0] aint_n[3] aint_n[4] aint_n[5] aint_n[6] DP8TDec_and4_x1
Xpage_and[1] vdd vss page[1] aint[3] aint_n[4] aint_n[5] aint_n[6] DP8TDec_and4_x1
Xpage_and[2] vdd vss page[2] aint_n[3] aint[4] aint_n[5] aint_n[6] DP8TDec_and4_x1
Xpage_and[3] vdd vss page[3] aint[3] aint[4] aint_n[5] aint_n[6] DP8TDec_and4_x1
Xpage_and[4] vdd vss page[4] aint_n[3] aint_n[4] aint[5] aint_n[6] DP8TDec_and4_x1
Xpage_and[5] vdd vss page[5] aint[3] aint_n[4] aint[5] aint_n[6] DP8TDec_and4_x1
Xpage_and[6] vdd vss page[6] aint_n[3] aint[4] aint[5] aint_n[6] DP8TDec_and4_x1
Xpage_and[7] vdd vss page[7] aint[3] aint[4] aint[5] aint_n[6] DP8TDec_and4_x1
Xpage_and[8] vdd vss page[8] aint_n[3] aint_n[4] aint_n[5] aint[6] DP8TDec_and4_x1
Xpage_and[9] vdd vss page[9] aint[3] aint_n[4] aint_n[5] aint[6] DP8TDec_and4_x1
Xpage_and[10] vdd vss page[10] aint_n[3] aint[4] aint_n[5] aint[6] DP8TDec_and4_x1
Xpage_and[11] vdd vss page[11] aint[3] aint[4] aint_n[5] aint[6] DP8TDec_and4_x1
Xpage_and[12] vdd vss page[12] aint_n[3] aint_n[4] aint[5] aint[6] DP8TDec_and4_x1
Xpage_and[13] vdd vss page[13] aint[3] aint_n[4] aint[5] aint[6] DP8TDec_and4_x1
Xpage_and[14] vdd vss page[14] aint_n[3] aint[4] aint[5] aint[6] DP8TDec_and4_x1
Xpage_and[15] vdd vss page[15] aint[3] aint[4] aint[5] aint[6] DP8TDec_and4_x1
.ends DP8TRowPredecoders_3_4B_wl2

.subckt DP8TWLDrive_26LN100WN26LP200WP_wl2 vss substrate vdd nwell wl_n wl_drive
Xnmos1 vss wl_n wl_drive substrate sg13_lv_nmos l=0.13um w=0.5um
Xnmos2 wl_drive wl_n vss substrate sg13_lv_nmos l=0.13um w=0.5um
Xpmos1 vdd wl_n wl_drive nwell sg13_lv_pmos l=0.13um w=1.0um
Xpmos2 wl_drive wl_n vdd nwell sg13_lv_pmos l=0.13um w=1.0um
.ends DP8TWLDrive_26LN100WN26LP200WP_wl2

.subckt DP8TRowDecoderDriverPage_2PD8R_wl2 vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page wl_en
Xnand3[0] vss vdd pd[0][0] pd[0][1] page wl_en wl_n[0] wl_n[1] DP8TRowDecoderNand3X2
Xnand3[1] vss vdd pd[0][2] pd[0][3] page wl_en wl_n[2] wl_n[3] DP8TRowDecoderNand3X2
Xnand3[2] vss vdd pd[0][4] pd[0][5] page wl_en wl_n[4] wl_n[5] DP8TRowDecoderNand3X2
Xnand3[3] vss vdd pd[0][6] pd[0][7] page wl_en wl_n[6] wl_n[7] DP8TRowDecoderNand3X2
Xdrive[0] vss vss vdd vdd wl_n[0] wl[0] DP8TWLDrive_26LN100WN26LP200WP_wl2
Xdrive[1] vss vss vdd vdd wl_n[1] wl[1] DP8TWLDrive_26LN100WN26LP200WP_wl2
Xdrive[2] vss vss vdd vdd wl_n[2] wl[2] DP8TWLDrive_26LN100WN26LP200WP_wl2
Xdrive[3] vss vss vdd vdd wl_n[3] wl[3] DP8TWLDrive_26LN100WN26LP200WP_wl2
Xdrive[4] vss vss vdd vdd wl_n[4] wl[4] DP8TWLDrive_26LN100WN26LP200WP_wl2
Xdrive[5] vss vss vdd vdd wl_n[5] wl[5] DP8TWLDrive_26LN100WN26LP200WP_wl2
Xdrive[6] vss vss vdd vdd wl_n[6] wl[6] DP8TWLDrive_26LN100WN26LP200WP_wl2
Xdrive[7] vss vss vdd vdd wl_n[7] wl[7] DP8TWLDrive_26LN100WN26LP200WP_wl2
.ends DP8TRowDecoderDriverPage_2PD8R_wl2

.subckt DP8TRowDecoder_3_4B_wl2 vss vdd a[0] a[1] a[2] a[3] a[4] a[5] a[6] clk wl_en wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127]
Xpredec vss vdd clk a[0] a[1] a[2] a[3] a[4] a[5] a[6] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[0] page[1] page[2] page[3] page[4] page[5] page[6] page[7] page[8] page[9] page[10] page[11] page[12] page[13] page[14] page[15] DP8TRowPredecoders_3_4B_wl2
Xpage[0] vss vdd wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[0] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[1] vss vdd wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[1] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[2] vss vdd wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[2] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[3] vss vdd wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[3] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[4] vss vdd wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[4] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[5] vss vdd wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[5] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[6] vss vdd wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[6] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[7] vss vdd wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[7] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[8] vss vdd wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[8] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[9] vss vdd wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[9] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[10] vss vdd wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[10] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[11] vss vdd wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[11] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[12] vss vdd wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[12] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[13] vss vdd wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[13] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[14] vss vdd wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[14] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xpage[15] vss vdd wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] pd[0][0] pd[0][1] pd[0][2] pd[0][3] pd[0][4] pd[0][5] pd[0][6] pd[0][7] page[15] wl_en DP8TRowDecoderDriverPage_2PD8R_wl2
Xbulkcon[0] vdd vss DP8TRowDecoderBulkConn
Xbulkcon[1] vdd vss DP8TRowDecoderBulkConn
Xbulkcon[2] vdd vss DP8TRowDecoderBulkConn
Xbulkcon[3] vdd vss DP8TRowDecoderBulkConn
Xbulkcon[4] vdd vss DP8TRowDecoderBulkConn
Xbulkcon[5] vdd vss DP8TRowDecoderBulkConn
Xbulkcon[6] vdd vss DP8TRowDecoderBulkConn
Xbulkcon[7] vdd vss DP8TRowDecoderBulkConn
Xbulkcon[8] vdd vss DP8TRowDecoderBulkConn
.ends DP8TRowDecoder_3_4B_wl2

.subckt DP8TRowPeriphery_3_4_2_wl2 vss vdd clk a[0] a[1] a[2] a[3] a[4] a[5] a[6] a[7] a[8] wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] mux[0] mux[1] mux[2] mux[3] columnclk precharge_n we_en
Xclkgen vss vdd clk decodeclk columnclk precharge_n wl_en we_en DP8TClockGenerator_8S1R
Xcoldec vss vdd decodeclk a[0] a[1] mux[0] mux[1] mux[2] mux[3] DP8TLatchedDecoder_2A2R
Xrowdec vss vdd a[2] a[3] a[4] a[5] a[6] a[7] a[8] decodeclk wl_en wl[0] wl[1] wl[2] wl[3] wl[4] wl[5] wl[6] wl[7] wl[8] wl[9] wl[10] wl[11] wl[12] wl[13] wl[14] wl[15] wl[16] wl[17] wl[18] wl[19] wl[20] wl[21] wl[22] wl[23] wl[24] wl[25] wl[26] wl[27] wl[28] wl[29] wl[30] wl[31] wl[32] wl[33] wl[34] wl[35] wl[36] wl[37] wl[38] wl[39] wl[40] wl[41] wl[42] wl[43] wl[44] wl[45] wl[46] wl[47] wl[48] wl[49] wl[50] wl[51] wl[52] wl[53] wl[54] wl[55] wl[56] wl[57] wl[58] wl[59] wl[60] wl[61] wl[62] wl[63] wl[64] wl[65] wl[66] wl[67] wl[68] wl[69] wl[70] wl[71] wl[72] wl[73] wl[74] wl[75] wl[76] wl[77] wl[78] wl[79] wl[80] wl[81] wl[82] wl[83] wl[84] wl[85] wl[86] wl[87] wl[88] wl[89] wl[90] wl[91] wl[92] wl[93] wl[94] wl[95] wl[96] wl[97] wl[98] wl[99] wl[100] wl[101] wl[102] wl[103] wl[104] wl[105] wl[106] wl[107] wl[108] wl[109] wl[110] wl[111] wl[112] wl[113] wl[114] wl[115] wl[116] wl[117] wl[118] wl[119] wl[120] wl[121] wl[122] wl[123] wl[124] wl[125] wl[126] wl[127] DP8TRowDecoder_3_4B_wl2
.ends DP8TRowPeriphery_3_4_2_wl2

.subckt DP8TCell vss substrate vdd nwell wl1 wl2 bl1 bl1_n bl2 bl2_n
Xpu1 vdd bit_n bit nwell sg13_lv_pmos l=0.13um w=0.15um
Xpd1 bit bit_n vss substrate sg13_lv_nmos l=0.13um w=0.2um
Xpu2 vdd bit bit_n nwell sg13_lv_pmos l=0.13um w=0.15um
Xpd2 bit_n bit vss substrate sg13_lv_nmos l=0.13um w=0.2um
Xpg1 bit wl1 bl1 substrate sg13_lv_nmos l=0.13um w=0.2um
Xpg1n bit_n wl1 bl1_n substrate sg13_lv_nmos l=0.13um w=0.2um
Xpg2 bit wl2 bl2 substrate sg13_lv_nmos l=0.13um w=0.2um
Xpg2n bit_n wl2 bl2_n substrate sg13_lv_nmos l=0.13um w=0.2um
.ends DP8TCell

.subckt DP8TArray_2X1 vss substrate vdd nwell wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0]
Xinst0x0 vss substrate vdd nwell wl1[0] wl2[0] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TCell
Xinst1x0 vss substrate vdd nwell wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TCell
.ends DP8TArray_2X1

.subckt DP8TArray_2X2 vss substrate vdd nwell wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss substrate vdd nwell wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] DP8TArray_2X1
Xinst0x1 vss substrate vdd nwell wl1[0] wl2[0] wl1[1] wl2[1] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TArray_2X1
.ends DP8TArray_2X2

.subckt DP8TArray_4X2 vss substrate vdd nwell wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0x0 vss substrate vdd nwell wl1[0] wl2[0] wl1[1] wl2[1] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TArray_2X2
Xinst1x0 vss substrate vdd nwell wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TArray_2X2
.ends DP8TArray_4X2

.subckt DP8TArray_4X4 vss substrate vdd nwell wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss substrate vdd nwell wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TArray_4X2
Xinst0x1 vss substrate vdd nwell wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TArray_4X2
.ends DP8TArray_4X4

.subckt DP8TArray_8X4 vss substrate vdd nwell wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0x0 vss substrate vdd nwell wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TArray_4X4
Xinst1x0 vss substrate vdd nwell wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TArray_4X4
.ends DP8TArray_8X4

.subckt DP8TArray_8X8 vss substrate vdd nwell wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss substrate vdd nwell wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TArray_8X4
Xinst0x1 vss substrate vdd nwell wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TArray_8X4
.ends DP8TArray_8X8

.subckt DP8TArray_16X8 vss substrate vdd nwell wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0x0 vss substrate vdd nwell wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TArray_8X8
Xinst1x0 vss substrate vdd nwell wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TArray_8X8
.ends DP8TArray_16X8

.subckt DP8TArray_16X16 vss substrate vdd nwell wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15]
Xinst0x0 vss substrate vdd nwell wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TArray_16X8
Xinst0x1 vss substrate vdd nwell wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] DP8TArray_16X8
.ends DP8TArray_16X16

.subckt DP8TArray_16X32 vss substrate vdd nwell wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31]
Xinst0x0 vss substrate vdd nwell wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] DP8TArray_16X16
Xinst0x1 vss substrate vdd nwell wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_16X16
.ends DP8TArray_16X32

.subckt DP8TBulkConnRow_32 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] DP8TBulkConnRow_16
Xinst1 vss vdd bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TBulkConnRow_16
.ends DP8TBulkConnRow_32

.subckt DP8TArray_32X32 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31]
Xinst0x0 vss vss vdd vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_16X32
Xinst1x0 vss vss vdd vdd wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_16X32
Xbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TBulkConnRow_32
.ends DP8TArray_32X32

.subckt DP8TArray_64X32 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_32X32
Xinst1x0 vss vdd wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_32X32
Xbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TBulkConnRow_32
.ends DP8TArray_64X32

.subckt DP8TBulkConn vdd vss bl1 bl2 bl1_n bl2_n

.ends DP8TBulkConn

.subckt DP8TBulkConnRow_2 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1]
Xinst0 vdd vss bl1[0] bl2[0] bl1_n[0] bl2_n[0] DP8TBulkConn
Xinst1 vdd vss bl1[1] bl2[1] bl1_n[1] bl2_n[1] DP8TBulkConn
.ends DP8TBulkConnRow_2

.subckt DP8TBulkConnRow_4 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] DP8TBulkConnRow_2
Xinst1 vss vdd bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TBulkConnRow_2
.ends DP8TBulkConnRow_4

.subckt DP8TBulkConnRow_8 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] DP8TBulkConnRow_4
Xinst1 vss vdd bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TBulkConnRow_4
.ends DP8TBulkConnRow_8

.subckt DP8TBulkConnRow_16 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15]
Xinst0 vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] DP8TBulkConnRow_8
Xinst1 vss vdd bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] DP8TBulkConnRow_8
.ends DP8TBulkConnRow_16

.subckt DP8TArray_128X32BC vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31]
Xinst0x0 vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_64X32
Xinst1x0 vss vdd wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_64X32
Xbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TBulkConnRow_32
Xbottombcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TBulkConnRow_32
Xtopbcrow vss vdd bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TBulkConnRow_32
.ends DP8TArray_128X32BC

.subckt DP8TPrecharge_bl1 vdd nwell bl bl_n precharge_n
Xpc1 vdd precharge_n bl nwell sg13_lv_pmos l=0.13um w=0.5um
Xpc2 bl precharge_n bl_n nwell sg13_lv_pmos l=0.13um w=0.5um
Xpc3 bl_n precharge_n vdd nwell sg13_lv_pmos l=0.13um w=0.5um
.ends DP8TPrecharge_bl1

.subckt DP8TColMux_4C26L699W_bl1 bl[0] bl_n[0] mux[0] bl[1] bl_n[1] mux[1] bl[2] bl_n[2] mux[2] bl[3] bl_n[3] mux[3] vss muxbl muxbl_n
Xpgbl0 muxbl mux[0] bl[0] vss sg13_lv_nmos l=0.13um w=3.5um
Xpgbln0 bl_n[0] mux[0] muxbl_n vss sg13_lv_nmos l=0.13um w=3.5um
Xpgbl1 bl[1] mux[1] muxbl vss sg13_lv_nmos l=0.13um w=3.5um
Xpgbln1 muxbl_n mux[1] bl_n[1] vss sg13_lv_nmos l=0.13um w=3.5um
Xpgbl2 muxbl mux[2] bl[2] vss sg13_lv_nmos l=0.13um w=3.5um
Xpgbln2 bl_n[2] mux[2] muxbl_n vss sg13_lv_nmos l=0.13um w=3.5um
Xpgbl3 bl[3] mux[3] muxbl vss sg13_lv_nmos l=0.13um w=3.5um
Xpgbln3 muxbl_n mux[3] bl_n[3] vss sg13_lv_nmos l=0.13um w=3.5um
.ends DP8TColMux_4C26L699W_bl1

.subckt DP8TReadWrite_4M vss vdd d q bl bl_n clk we_n
Xsenseamp vdd vss bl_n bl q noconn nsnrlatch_x1
Xd_ff vdd vss d clk d_l dff_x1
Xd_inv vdd vss d_l d_n inv_x0
Xnora vdd vss bl_pd_g d_l we_n nor2_x0
Xnorb vdd vss bln_pd_g d_n we_n nor2_x0
Xbl_pd bl bl_pd_g vss vss sg13_lv_nmos l=0.13um w=1.9um
Xbln_pd vss bln_pd_g bl_n vss sg13_lv_nmos l=0.13um w=1.9um
.ends DP8TReadWrite_4M

.subckt DP8TClockWE vss vdd clkup clkdown we we_en we_n
Xclkbuf vdd vss clkup clkdown buf_x2
Xweff vdd vss we clkdown we_l dff_x1
Xwenand vdd vss we_n we_l we_en nand2_x0
.ends DP8TClockWE

.subckt DP8TColumnPeriphery_8B4M_bl1 vss vdd nwell clk precharge_n we we_en q[0] d[0] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] q[1] d[1] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] q[2] d[2] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] q[3] d[3] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15] q[4] d[4] bl[16] bl_n[16] bl[17] bl_n[17] bl[18] bl_n[18] bl[19] bl_n[19] q[5] d[5] bl[20] bl_n[20] bl[21] bl_n[21] bl[22] bl_n[22] bl[23] bl_n[23] q[6] d[6] bl[24] bl_n[24] bl[25] bl_n[25] bl[26] bl_n[26] bl[27] bl_n[27] q[7] d[7] bl[28] bl_n[28] bl[29] bl_n[29] bl[30] bl_n[30] bl[31] bl_n[31] mux[0] mux[1] mux[2] mux[3]
Xprecharge[0] vdd nwell bl[0] bl_n[0] precharge_n DP8TPrecharge_bl1
Xprecharge[1] vdd nwell bl[1] bl_n[1] precharge_n DP8TPrecharge_bl1
Xprecharge[2] vdd nwell bl[2] bl_n[2] precharge_n DP8TPrecharge_bl1
Xprecharge[3] vdd nwell bl[3] bl_n[3] precharge_n DP8TPrecharge_bl1
Xprecharge[4] vdd nwell bl[4] bl_n[4] precharge_n DP8TPrecharge_bl1
Xprecharge[5] vdd nwell bl[5] bl_n[5] precharge_n DP8TPrecharge_bl1
Xprecharge[6] vdd nwell bl[6] bl_n[6] precharge_n DP8TPrecharge_bl1
Xprecharge[7] vdd nwell bl[7] bl_n[7] precharge_n DP8TPrecharge_bl1
Xprecharge[8] vdd nwell bl[8] bl_n[8] precharge_n DP8TPrecharge_bl1
Xprecharge[9] vdd nwell bl[9] bl_n[9] precharge_n DP8TPrecharge_bl1
Xprecharge[10] vdd nwell bl[10] bl_n[10] precharge_n DP8TPrecharge_bl1
Xprecharge[11] vdd nwell bl[11] bl_n[11] precharge_n DP8TPrecharge_bl1
Xprecharge[12] vdd nwell bl[12] bl_n[12] precharge_n DP8TPrecharge_bl1
Xprecharge[13] vdd nwell bl[13] bl_n[13] precharge_n DP8TPrecharge_bl1
Xprecharge[14] vdd nwell bl[14] bl_n[14] precharge_n DP8TPrecharge_bl1
Xprecharge[15] vdd nwell bl[15] bl_n[15] precharge_n DP8TPrecharge_bl1
Xprecharge[16] vdd nwell bl[16] bl_n[16] precharge_n DP8TPrecharge_bl1
Xprecharge[17] vdd nwell bl[17] bl_n[17] precharge_n DP8TPrecharge_bl1
Xprecharge[18] vdd nwell bl[18] bl_n[18] precharge_n DP8TPrecharge_bl1
Xprecharge[19] vdd nwell bl[19] bl_n[19] precharge_n DP8TPrecharge_bl1
Xprecharge[20] vdd nwell bl[20] bl_n[20] precharge_n DP8TPrecharge_bl1
Xprecharge[21] vdd nwell bl[21] bl_n[21] precharge_n DP8TPrecharge_bl1
Xprecharge[22] vdd nwell bl[22] bl_n[22] precharge_n DP8TPrecharge_bl1
Xprecharge[23] vdd nwell bl[23] bl_n[23] precharge_n DP8TPrecharge_bl1
Xprecharge[24] vdd nwell bl[24] bl_n[24] precharge_n DP8TPrecharge_bl1
Xprecharge[25] vdd nwell bl[25] bl_n[25] precharge_n DP8TPrecharge_bl1
Xprecharge[26] vdd nwell bl[26] bl_n[26] precharge_n DP8TPrecharge_bl1
Xprecharge[27] vdd nwell bl[27] bl_n[27] precharge_n DP8TPrecharge_bl1
Xprecharge[28] vdd nwell bl[28] bl_n[28] precharge_n DP8TPrecharge_bl1
Xprecharge[29] vdd nwell bl[29] bl_n[29] precharge_n DP8TPrecharge_bl1
Xprecharge[30] vdd nwell bl[30] bl_n[30] precharge_n DP8TPrecharge_bl1
Xprecharge[31] vdd nwell bl[31] bl_n[31] precharge_n DP8TPrecharge_bl1
Xcolmux[0] bl[0] bl_n[0] mux[0] bl[1] bl_n[1] mux[1] bl[2] bl_n[2] mux[2] bl[3] bl_n[3] mux[3] vss muxbl[0] muxbl_n[0] DP8TColMux_4C26L699W_bl1
Xcolmux[1] bl[4] bl_n[4] mux[0] bl[5] bl_n[5] mux[1] bl[6] bl_n[6] mux[2] bl[7] bl_n[7] mux[3] vss muxbl[1] muxbl_n[1] DP8TColMux_4C26L699W_bl1
Xcolmux[2] bl[8] bl_n[8] mux[0] bl[9] bl_n[9] mux[1] bl[10] bl_n[10] mux[2] bl[11] bl_n[11] mux[3] vss muxbl[2] muxbl_n[2] DP8TColMux_4C26L699W_bl1
Xcolmux[3] bl[12] bl_n[12] mux[0] bl[13] bl_n[13] mux[1] bl[14] bl_n[14] mux[2] bl[15] bl_n[15] mux[3] vss muxbl[3] muxbl_n[3] DP8TColMux_4C26L699W_bl1
Xcolmux[4] bl[16] bl_n[16] mux[0] bl[17] bl_n[17] mux[1] bl[18] bl_n[18] mux[2] bl[19] bl_n[19] mux[3] vss muxbl[4] muxbl_n[4] DP8TColMux_4C26L699W_bl1
Xcolmux[5] bl[20] bl_n[20] mux[0] bl[21] bl_n[21] mux[1] bl[22] bl_n[22] mux[2] bl[23] bl_n[23] mux[3] vss muxbl[5] muxbl_n[5] DP8TColMux_4C26L699W_bl1
Xcolmux[6] bl[24] bl_n[24] mux[0] bl[25] bl_n[25] mux[1] bl[26] bl_n[26] mux[2] bl[27] bl_n[27] mux[3] vss muxbl[6] muxbl_n[6] DP8TColMux_4C26L699W_bl1
Xcolmux[7] bl[28] bl_n[28] mux[0] bl[29] bl_n[29] mux[1] bl[30] bl_n[30] mux[2] bl[31] bl_n[31] mux[3] vss muxbl[7] muxbl_n[7] DP8TColMux_4C26L699W_bl1
Xrw[0] vss vdd d[0] q[0] muxbl[0] muxbl_n[0] intclk we_n DP8TReadWrite_4M
Xrw[1] vss vdd d[1] q[1] muxbl[1] muxbl_n[1] intclk we_n DP8TReadWrite_4M
Xrw[2] vss vdd d[2] q[2] muxbl[2] muxbl_n[2] intclk we_n DP8TReadWrite_4M
Xrw[3] vss vdd d[3] q[3] muxbl[3] muxbl_n[3] intclk we_n DP8TReadWrite_4M
Xrw[4] vss vdd d[4] q[4] muxbl[4] muxbl_n[4] intclk we_n DP8TReadWrite_4M
Xrw[5] vss vdd d[5] q[5] muxbl[5] muxbl_n[5] intclk we_n DP8TReadWrite_4M
Xrw[6] vss vdd d[6] q[6] muxbl[6] muxbl_n[6] intclk we_n DP8TReadWrite_4M
Xrw[7] vss vdd d[7] q[7] muxbl[7] muxbl_n[7] intclk we_n DP8TReadWrite_4M
Xclkwe vss vdd clk intclk we we_en we_n DP8TClockWE
.ends DP8TColumnPeriphery_8B4M_bl1

.subckt DP8TPrecharge_bl2 vdd nwell bl bl_n precharge_n
Xpc1 vdd precharge_n bl nwell sg13_lv_pmos l=0.13um w=0.5um
Xpc2 bl precharge_n bl_n nwell sg13_lv_pmos l=0.13um w=0.5um
Xpc3 bl_n precharge_n vdd nwell sg13_lv_pmos l=0.13um w=0.5um
.ends DP8TPrecharge_bl2

.subckt DP8TColMux_4C26L699WR_bl2 bl[3] bl_n[3] mux[3] bl[2] bl_n[2] mux[2] bl[1] bl_n[1] mux[1] bl[0] bl_n[0] mux[0] vss muxbl muxbl_n
Xpgbl3 muxbl mux[3] bl[3] vss sg13_lv_nmos l=0.13um w=3.5um
Xpgbln3 bl_n[3] mux[3] muxbl_n vss sg13_lv_nmos l=0.13um w=3.5um
Xpgbl2 bl[2] mux[2] muxbl vss sg13_lv_nmos l=0.13um w=3.5um
Xpgbln2 muxbl_n mux[2] bl_n[2] vss sg13_lv_nmos l=0.13um w=3.5um
Xpgbl1 muxbl mux[1] bl[1] vss sg13_lv_nmos l=0.13um w=3.5um
Xpgbln1 bl_n[1] mux[1] muxbl_n vss sg13_lv_nmos l=0.13um w=3.5um
Xpgbl0 bl[0] mux[0] muxbl vss sg13_lv_nmos l=0.13um w=3.5um
Xpgbln0 muxbl_n mux[0] bl_n[0] vss sg13_lv_nmos l=0.13um w=3.5um
.ends DP8TColMux_4C26L699WR_bl2

.subckt nsnrlatch_x1 vdd vss nset nrst q nq
Xnset_nmos q nset _net0 vss sg13_lv_nmos l=0.13um w=1.31um
Xnset_pmos vdd nset q vdd sg13_lv_pmos l=0.13um w=1.3um
Xnq_nmos _net0 nq vss vss sg13_lv_nmos l=0.13um w=1.31um
Xnq_pmos q nq vdd vdd sg13_lv_pmos l=0.13um w=1.3um
Xq_nmos vss q _net1 vss sg13_lv_nmos l=0.13um w=1.31um
Xq_pmos vdd q nq vdd sg13_lv_pmos l=0.13um w=1.3um
Xnrst_nmos _net1 nrst nq vss sg13_lv_nmos l=0.13um w=1.31um
Xnrst_pmos nq nrst vdd vdd sg13_lv_pmos l=0.13um w=1.3um
.ends nsnrlatch_x1

.subckt dff_x1 vdd vss i clk q
Xclk_nmos _clk_n clk vss vss sg13_lv_nmos l=0.13um w=0.78um
Xclk_pmos _clk_n clk vdd vdd sg13_lv_pmos l=0.13um w=0.78um
Xclk_n_nmos0 vss _clk_n _clk_buf vss sg13_lv_nmos l=0.13um w=0.78um
Xclk_n_pmos0 vdd _clk_n _clk_buf vdd sg13_lv_pmos l=0.13um w=0.78um
Xi_nmos _u i vss vss sg13_lv_nmos l=0.13um w=0.78um
Xi_pmos _u i vdd vdd sg13_lv_pmos l=0.13um w=0.78um
Xu_nmos vss _u _net0 vss sg13_lv_nmos l=0.13um w=0.78um
Xu_pmos vdd _u _net1 vdd sg13_lv_pmos l=0.13um w=0.78um
Xclk_n_nmos1 _net0 _clk_n _dff_m vss sg13_lv_nmos l=0.13um w=0.78um
Xclk_buf_pmos0 _net1 _clk_buf _dff_m vdd sg13_lv_pmos l=0.13um w=0.78um
Xclk_buf_nmos0 _dff_m _clk_buf _net2 vss sg13_lv_nmos l=0.13um w=0.78um
Xclk_n_pmos1 _dff_m _clk_n _net3 vdd sg13_lv_pmos l=0.13um w=0.78um
Xy_nmos _net2 _y vss vss sg13_lv_nmos l=0.13um w=0.78um
Xy_pmos _net3 _y vdd vdd sg13_lv_pmos l=0.13um w=0.78um
Xdff_m_nmos vss _dff_m _y vss sg13_lv_nmos l=0.13um w=0.78um
Xdff_m_pmos vdd _dff_m _y vdd sg13_lv_pmos l=0.13um w=0.78um
Xclk_buf_nmos1 _y _clk_buf _dff_s vss sg13_lv_nmos l=0.13um w=0.78um
Xclk_n_pmos2 _y _clk_n _dff_s vdd sg13_lv_pmos l=0.13um w=0.78um
Xclk_n_nmos2 _dff_s _clk_n _net4 vss sg13_lv_nmos l=0.13um w=0.78um
Xclk_buf_pmos1 _dff_s _clk_buf _net5 vdd sg13_lv_pmos l=0.13um w=0.78um
Xq_nmos _net4 q vss vss sg13_lv_nmos l=0.13um w=0.78um
Xq_pmos _net5 q vdd vdd sg13_lv_pmos l=0.13um w=0.78um
Xdff_s_nmos vss _dff_s q vss sg13_lv_nmos l=0.13um w=0.83um
Xdff_s_pmos vdd _dff_s q vdd sg13_lv_pmos l=0.13um w=0.82um
.ends dff_x1

.subckt nor2_x0 vdd vss nq i0 i1
Xi0_nmos vss i0 nq vss sg13_lv_nmos l=0.13um w=0.78um
Xi0_pmos vdd i0 _net0 vdd sg13_lv_pmos l=0.13um w=0.78um
Xi1_nmos nq i1 vss vss sg13_lv_nmos l=0.13um w=0.78um
Xi1_pmos _net0 i1 nq vdd sg13_lv_pmos l=0.13um w=0.78um
.ends nor2_x0

.subckt buf_x2 vdd vss i q
Xstage0_nmos _i_n i vss vss sg13_lv_nmos l=0.13um w=0.78um
Xstage0_pmos _i_n i vdd vdd sg13_lv_pmos l=0.13um w=0.78um
Xnmos[0] vss _i_n q vss sg13_lv_nmos l=0.13um w=1.07um
Xpmos[0] vdd _i_n q vdd sg13_lv_pmos l=0.13um w=1.06um
Xnmos[1] q _i_n vss vss sg13_lv_nmos l=0.13um w=1.07um
Xpmos[1] q _i_n vdd vdd sg13_lv_pmos l=0.13um w=1.06um
.ends buf_x2

.subckt DP8TColumnPeriphery_8B4MR_bl2 vss vdd nwell clk precharge_n we we_en q[0] d[0] bl[0] bl_n[0] bl[1] bl_n[1] bl[2] bl_n[2] bl[3] bl_n[3] q[1] d[1] bl[4] bl_n[4] bl[5] bl_n[5] bl[6] bl_n[6] bl[7] bl_n[7] q[2] d[2] bl[8] bl_n[8] bl[9] bl_n[9] bl[10] bl_n[10] bl[11] bl_n[11] q[3] d[3] bl[12] bl_n[12] bl[13] bl_n[13] bl[14] bl_n[14] bl[15] bl_n[15] q[4] d[4] bl[16] bl_n[16] bl[17] bl_n[17] bl[18] bl_n[18] bl[19] bl_n[19] q[5] d[5] bl[20] bl_n[20] bl[21] bl_n[21] bl[22] bl_n[22] bl[23] bl_n[23] q[6] d[6] bl[24] bl_n[24] bl[25] bl_n[25] bl[26] bl_n[26] bl[27] bl_n[27] q[7] d[7] bl[28] bl_n[28] bl[29] bl_n[29] bl[30] bl_n[30] bl[31] bl_n[31] mux[0] mux[1] mux[2] mux[3]
Xprecharge[0] vdd nwell bl[0] bl_n[0] precharge_n DP8TPrecharge_bl2
Xprecharge[1] vdd nwell bl[1] bl_n[1] precharge_n DP8TPrecharge_bl2
Xprecharge[2] vdd nwell bl[2] bl_n[2] precharge_n DP8TPrecharge_bl2
Xprecharge[3] vdd nwell bl[3] bl_n[3] precharge_n DP8TPrecharge_bl2
Xprecharge[4] vdd nwell bl[4] bl_n[4] precharge_n DP8TPrecharge_bl2
Xprecharge[5] vdd nwell bl[5] bl_n[5] precharge_n DP8TPrecharge_bl2
Xprecharge[6] vdd nwell bl[6] bl_n[6] precharge_n DP8TPrecharge_bl2
Xprecharge[7] vdd nwell bl[7] bl_n[7] precharge_n DP8TPrecharge_bl2
Xprecharge[8] vdd nwell bl[8] bl_n[8] precharge_n DP8TPrecharge_bl2
Xprecharge[9] vdd nwell bl[9] bl_n[9] precharge_n DP8TPrecharge_bl2
Xprecharge[10] vdd nwell bl[10] bl_n[10] precharge_n DP8TPrecharge_bl2
Xprecharge[11] vdd nwell bl[11] bl_n[11] precharge_n DP8TPrecharge_bl2
Xprecharge[12] vdd nwell bl[12] bl_n[12] precharge_n DP8TPrecharge_bl2
Xprecharge[13] vdd nwell bl[13] bl_n[13] precharge_n DP8TPrecharge_bl2
Xprecharge[14] vdd nwell bl[14] bl_n[14] precharge_n DP8TPrecharge_bl2
Xprecharge[15] vdd nwell bl[15] bl_n[15] precharge_n DP8TPrecharge_bl2
Xprecharge[16] vdd nwell bl[16] bl_n[16] precharge_n DP8TPrecharge_bl2
Xprecharge[17] vdd nwell bl[17] bl_n[17] precharge_n DP8TPrecharge_bl2
Xprecharge[18] vdd nwell bl[18] bl_n[18] precharge_n DP8TPrecharge_bl2
Xprecharge[19] vdd nwell bl[19] bl_n[19] precharge_n DP8TPrecharge_bl2
Xprecharge[20] vdd nwell bl[20] bl_n[20] precharge_n DP8TPrecharge_bl2
Xprecharge[21] vdd nwell bl[21] bl_n[21] precharge_n DP8TPrecharge_bl2
Xprecharge[22] vdd nwell bl[22] bl_n[22] precharge_n DP8TPrecharge_bl2
Xprecharge[23] vdd nwell bl[23] bl_n[23] precharge_n DP8TPrecharge_bl2
Xprecharge[24] vdd nwell bl[24] bl_n[24] precharge_n DP8TPrecharge_bl2
Xprecharge[25] vdd nwell bl[25] bl_n[25] precharge_n DP8TPrecharge_bl2
Xprecharge[26] vdd nwell bl[26] bl_n[26] precharge_n DP8TPrecharge_bl2
Xprecharge[27] vdd nwell bl[27] bl_n[27] precharge_n DP8TPrecharge_bl2
Xprecharge[28] vdd nwell bl[28] bl_n[28] precharge_n DP8TPrecharge_bl2
Xprecharge[29] vdd nwell bl[29] bl_n[29] precharge_n DP8TPrecharge_bl2
Xprecharge[30] vdd nwell bl[30] bl_n[30] precharge_n DP8TPrecharge_bl2
Xprecharge[31] vdd nwell bl[31] bl_n[31] precharge_n DP8TPrecharge_bl2
Xcolmux[0] bl[3] bl_n[3] mux[3] bl[2] bl_n[2] mux[2] bl[1] bl_n[1] mux[1] bl[0] bl_n[0] mux[0] vss muxbl[0] muxbl_n[0] DP8TColMux_4C26L699WR_bl2
Xcolmux[1] bl[7] bl_n[7] mux[3] bl[6] bl_n[6] mux[2] bl[5] bl_n[5] mux[1] bl[4] bl_n[4] mux[0] vss muxbl[1] muxbl_n[1] DP8TColMux_4C26L699WR_bl2
Xcolmux[2] bl[11] bl_n[11] mux[3] bl[10] bl_n[10] mux[2] bl[9] bl_n[9] mux[1] bl[8] bl_n[8] mux[0] vss muxbl[2] muxbl_n[2] DP8TColMux_4C26L699WR_bl2
Xcolmux[3] bl[15] bl_n[15] mux[3] bl[14] bl_n[14] mux[2] bl[13] bl_n[13] mux[1] bl[12] bl_n[12] mux[0] vss muxbl[3] muxbl_n[3] DP8TColMux_4C26L699WR_bl2
Xcolmux[4] bl[19] bl_n[19] mux[3] bl[18] bl_n[18] mux[2] bl[17] bl_n[17] mux[1] bl[16] bl_n[16] mux[0] vss muxbl[4] muxbl_n[4] DP8TColMux_4C26L699WR_bl2
Xcolmux[5] bl[23] bl_n[23] mux[3] bl[22] bl_n[22] mux[2] bl[21] bl_n[21] mux[1] bl[20] bl_n[20] mux[0] vss muxbl[5] muxbl_n[5] DP8TColMux_4C26L699WR_bl2
Xcolmux[6] bl[27] bl_n[27] mux[3] bl[26] bl_n[26] mux[2] bl[25] bl_n[25] mux[1] bl[24] bl_n[24] mux[0] vss muxbl[6] muxbl_n[6] DP8TColMux_4C26L699WR_bl2
Xcolmux[7] bl[31] bl_n[31] mux[3] bl[30] bl_n[30] mux[2] bl[29] bl_n[29] mux[1] bl[28] bl_n[28] mux[0] vss muxbl[7] muxbl_n[7] DP8TColMux_4C26L699WR_bl2
Xrw[0] vss vdd d[0] q[0] muxbl[0] muxbl_n[0] intclk we_n DP8TReadWrite_4M
Xrw[1] vss vdd d[1] q[1] muxbl[1] muxbl_n[1] intclk we_n DP8TReadWrite_4M
Xrw[2] vss vdd d[2] q[2] muxbl[2] muxbl_n[2] intclk we_n DP8TReadWrite_4M
Xrw[3] vss vdd d[3] q[3] muxbl[3] muxbl_n[3] intclk we_n DP8TReadWrite_4M
Xrw[4] vss vdd d[4] q[4] muxbl[4] muxbl_n[4] intclk we_n DP8TReadWrite_4M
Xrw[5] vss vdd d[5] q[5] muxbl[5] muxbl_n[5] intclk we_n DP8TReadWrite_4M
Xrw[6] vss vdd d[6] q[6] muxbl[6] muxbl_n[6] intclk we_n DP8TReadWrite_4M
Xrw[7] vss vdd d[7] q[7] muxbl[7] muxbl_n[7] intclk we_n DP8TReadWrite_4M
Xclkwe vss vdd clk intclk we we_en we_n DP8TClockWE
.ends DP8TColumnPeriphery_8B4MR_bl2

.subckt DP8TColumn_128R8B4M vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] q1[0] q2[0] d1[0] d2[0] q1[1] q2[1] d1[1] d2[1] q1[2] q2[2] d1[2] d2[2] q1[3] q2[3] d1[3] d2[3] q1[4] q2[4] d1[4] d2[4] q1[5] q2[5] d1[5] d2[5] q1[6] q2[6] d1[6] d2[6] q1[7] q2[7] d1[7] d2[7] we1 clk1 we_en1 precharge1_n we2 clk2 we_en2 precharge2_n mux1[0] mux2[0] mux1[1] mux2[1] mux1[2] mux2[2] mux1[3] mux2[3]
Xarray vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] bl1[0] bl1_n[0] bl2[0] bl2_n[0] bl1[1] bl1_n[1] bl2[1] bl2_n[1] bl1[2] bl1_n[2] bl2[2] bl2_n[2] bl1[3] bl1_n[3] bl2[3] bl2_n[3] bl1[4] bl1_n[4] bl2[4] bl2_n[4] bl1[5] bl1_n[5] bl2[5] bl2_n[5] bl1[6] bl1_n[6] bl2[6] bl2_n[6] bl1[7] bl1_n[7] bl2[7] bl2_n[7] bl1[8] bl1_n[8] bl2[8] bl2_n[8] bl1[9] bl1_n[9] bl2[9] bl2_n[9] bl1[10] bl1_n[10] bl2[10] bl2_n[10] bl1[11] bl1_n[11] bl2[11] bl2_n[11] bl1[12] bl1_n[12] bl2[12] bl2_n[12] bl1[13] bl1_n[13] bl2[13] bl2_n[13] bl1[14] bl1_n[14] bl2[14] bl2_n[14] bl1[15] bl1_n[15] bl2[15] bl2_n[15] bl1[16] bl1_n[16] bl2[16] bl2_n[16] bl1[17] bl1_n[17] bl2[17] bl2_n[17] bl1[18] bl1_n[18] bl2[18] bl2_n[18] bl1[19] bl1_n[19] bl2[19] bl2_n[19] bl1[20] bl1_n[20] bl2[20] bl2_n[20] bl1[21] bl1_n[21] bl2[21] bl2_n[21] bl1[22] bl1_n[22] bl2[22] bl2_n[22] bl1[23] bl1_n[23] bl2[23] bl2_n[23] bl1[24] bl1_n[24] bl2[24] bl2_n[24] bl1[25] bl1_n[25] bl2[25] bl2_n[25] bl1[26] bl1_n[26] bl2[26] bl2_n[26] bl1[27] bl1_n[27] bl2[27] bl2_n[27] bl1[28] bl1_n[28] bl2[28] bl2_n[28] bl1[29] bl1_n[29] bl2[29] bl2_n[29] bl1[30] bl1_n[30] bl2[30] bl2_n[30] bl1[31] bl1_n[31] bl2[31] bl2_n[31] DP8TArray_128X32BC
Xperiph1 vss vdd vdd clk1 precharge1_n we1 we_en1 q1[0] d1[0] bl1[0] bl1_n[0] bl1[1] bl1_n[1] bl1[2] bl1_n[2] bl1[3] bl1_n[3] q1[1] d1[1] bl1[4] bl1_n[4] bl1[5] bl1_n[5] bl1[6] bl1_n[6] bl1[7] bl1_n[7] q1[2] d1[2] bl1[8] bl1_n[8] bl1[9] bl1_n[9] bl1[10] bl1_n[10] bl1[11] bl1_n[11] q1[3] d1[3] bl1[12] bl1_n[12] bl1[13] bl1_n[13] bl1[14] bl1_n[14] bl1[15] bl1_n[15] q1[4] d1[4] bl1[16] bl1_n[16] bl1[17] bl1_n[17] bl1[18] bl1_n[18] bl1[19] bl1_n[19] q1[5] d1[5] bl1[20] bl1_n[20] bl1[21] bl1_n[21] bl1[22] bl1_n[22] bl1[23] bl1_n[23] q1[6] d1[6] bl1[24] bl1_n[24] bl1[25] bl1_n[25] bl1[26] bl1_n[26] bl1[27] bl1_n[27] q1[7] d1[7] bl1[28] bl1_n[28] bl1[29] bl1_n[29] bl1[30] bl1_n[30] bl1[31] bl1_n[31] mux1[0] mux1[1] mux1[2] mux1[3] DP8TColumnPeriphery_8B4M_bl1
Xperiph2 vss vdd vdd clk2 precharge2_n we2 we_en2 q2[0] d2[0] bl2[0] bl2_n[0] bl2[1] bl2_n[1] bl2[2] bl2_n[2] bl2[3] bl2_n[3] q2[1] d2[1] bl2[4] bl2_n[4] bl2[5] bl2_n[5] bl2[6] bl2_n[6] bl2[7] bl2_n[7] q2[2] d2[2] bl2[8] bl2_n[8] bl2[9] bl2_n[9] bl2[10] bl2_n[10] bl2[11] bl2_n[11] q2[3] d2[3] bl2[12] bl2_n[12] bl2[13] bl2_n[13] bl2[14] bl2_n[14] bl2[15] bl2_n[15] q2[4] d2[4] bl2[16] bl2_n[16] bl2[17] bl2_n[17] bl2[18] bl2_n[18] bl2[19] bl2_n[19] q2[5] d2[5] bl2[20] bl2_n[20] bl2[21] bl2_n[21] bl2[22] bl2_n[22] bl2[23] bl2_n[23] q2[6] d2[6] bl2[24] bl2_n[24] bl2[25] bl2_n[25] bl2[26] bl2_n[26] bl2[27] bl2_n[27] q2[7] d2[7] bl2[28] bl2_n[28] bl2[29] bl2_n[29] bl2[30] bl2_n[30] bl2[31] bl2_n[31] mux2[0] mux2[1] mux2[2] mux2[3] DP8TColumnPeriphery_8B4MR_bl2
.ends DP8TColumn_128R8B4M

.subckt DP8TColumnBlock_128R8B4M1W vss vdd clk1 clk2 precharge1_n precharge2_n we_en1 we_en2 wl1[0] wl1[1] wl1[2] wl1[3] wl1[4] wl1[5] wl1[6] wl1[7] wl1[8] wl1[9] wl1[10] wl1[11] wl1[12] wl1[13] wl1[14] wl1[15] wl1[16] wl1[17] wl1[18] wl1[19] wl1[20] wl1[21] wl1[22] wl1[23] wl1[24] wl1[25] wl1[26] wl1[27] wl1[28] wl1[29] wl1[30] wl1[31] wl1[32] wl1[33] wl1[34] wl1[35] wl1[36] wl1[37] wl1[38] wl1[39] wl1[40] wl1[41] wl1[42] wl1[43] wl1[44] wl1[45] wl1[46] wl1[47] wl1[48] wl1[49] wl1[50] wl1[51] wl1[52] wl1[53] wl1[54] wl1[55] wl1[56] wl1[57] wl1[58] wl1[59] wl1[60] wl1[61] wl1[62] wl1[63] wl1[64] wl1[65] wl1[66] wl1[67] wl1[68] wl1[69] wl1[70] wl1[71] wl1[72] wl1[73] wl1[74] wl1[75] wl1[76] wl1[77] wl1[78] wl1[79] wl1[80] wl1[81] wl1[82] wl1[83] wl1[84] wl1[85] wl1[86] wl1[87] wl1[88] wl1[89] wl1[90] wl1[91] wl1[92] wl1[93] wl1[94] wl1[95] wl1[96] wl1[97] wl1[98] wl1[99] wl1[100] wl1[101] wl1[102] wl1[103] wl1[104] wl1[105] wl1[106] wl1[107] wl1[108] wl1[109] wl1[110] wl1[111] wl1[112] wl1[113] wl1[114] wl1[115] wl1[116] wl1[117] wl1[118] wl1[119] wl1[120] wl1[121] wl1[122] wl1[123] wl1[124] wl1[125] wl1[126] wl1[127] wl2[0] wl2[1] wl2[2] wl2[3] wl2[4] wl2[5] wl2[6] wl2[7] wl2[8] wl2[9] wl2[10] wl2[11] wl2[12] wl2[13] wl2[14] wl2[15] wl2[16] wl2[17] wl2[18] wl2[19] wl2[20] wl2[21] wl2[22] wl2[23] wl2[24] wl2[25] wl2[26] wl2[27] wl2[28] wl2[29] wl2[30] wl2[31] wl2[32] wl2[33] wl2[34] wl2[35] wl2[36] wl2[37] wl2[38] wl2[39] wl2[40] wl2[41] wl2[42] wl2[43] wl2[44] wl2[45] wl2[46] wl2[47] wl2[48] wl2[49] wl2[50] wl2[51] wl2[52] wl2[53] wl2[54] wl2[55] wl2[56] wl2[57] wl2[58] wl2[59] wl2[60] wl2[61] wl2[62] wl2[63] wl2[64] wl2[65] wl2[66] wl2[67] wl2[68] wl2[69] wl2[70] wl2[71] wl2[72] wl2[73] wl2[74] wl2[75] wl2[76] wl2[77] wl2[78] wl2[79] wl2[80] wl2[81] wl2[82] wl2[83] wl2[84] wl2[85] wl2[86] wl2[87] wl2[88] wl2[89] wl2[90] wl2[91] wl2[92] wl2[93] wl2[94] wl2[95] wl2[96] wl2[97] wl2[98] wl2[99] wl2[100] wl2[101] wl2[102] wl2[103] wl2[104] wl2[105] wl2[106] wl2[107] wl2[108] wl2[109] wl2[110] wl2[111] wl2[112] wl2[113] wl2[114] wl2[115] wl2[116] wl2[117] wl2[118] wl2[119] wl2[120] wl2[121] wl2[122] wl2[123] wl2[124] wl2[125] wl2[126] wl2[127] mux1[0] mux1[1] mux1[2] mux1[3] mux2[0] mux2[1] mux2[2] mux2[3] we1[0] we2[0] q1[0] q2[0] d1[0] d2[0] q1[1] q2[1] d1[1] d2[1] q1[2] q2[2] d1[2] d2[2] q1[3] q2[3] d1[3] d2[3] q1[4] q2[4] d1[4] d2[4] q1[5] q2[5] d1[5] d2[5] q1[6] q2[6] d1[6] d2[6] q1[7] q2[7] d1[7] d2[7]
Xcolumn[0] vss vdd wl1[0] wl2[0] wl1[1] wl2[1] wl1[2] wl2[2] wl1[3] wl2[3] wl1[4] wl2[4] wl1[5] wl2[5] wl1[6] wl2[6] wl1[7] wl2[7] wl1[8] wl2[8] wl1[9] wl2[9] wl1[10] wl2[10] wl1[11] wl2[11] wl1[12] wl2[12] wl1[13] wl2[13] wl1[14] wl2[14] wl1[15] wl2[15] wl1[16] wl2[16] wl1[17] wl2[17] wl1[18] wl2[18] wl1[19] wl2[19] wl1[20] wl2[20] wl1[21] wl2[21] wl1[22] wl2[22] wl1[23] wl2[23] wl1[24] wl2[24] wl1[25] wl2[25] wl1[26] wl2[26] wl1[27] wl2[27] wl1[28] wl2[28] wl1[29] wl2[29] wl1[30] wl2[30] wl1[31] wl2[31] wl1[32] wl2[32] wl1[33] wl2[33] wl1[34] wl2[34] wl1[35] wl2[35] wl1[36] wl2[36] wl1[37] wl2[37] wl1[38] wl2[38] wl1[39] wl2[39] wl1[40] wl2[40] wl1[41] wl2[41] wl1[42] wl2[42] wl1[43] wl2[43] wl1[44] wl2[44] wl1[45] wl2[45] wl1[46] wl2[46] wl1[47] wl2[47] wl1[48] wl2[48] wl1[49] wl2[49] wl1[50] wl2[50] wl1[51] wl2[51] wl1[52] wl2[52] wl1[53] wl2[53] wl1[54] wl2[54] wl1[55] wl2[55] wl1[56] wl2[56] wl1[57] wl2[57] wl1[58] wl2[58] wl1[59] wl2[59] wl1[60] wl2[60] wl1[61] wl2[61] wl1[62] wl2[62] wl1[63] wl2[63] wl1[64] wl2[64] wl1[65] wl2[65] wl1[66] wl2[66] wl1[67] wl2[67] wl1[68] wl2[68] wl1[69] wl2[69] wl1[70] wl2[70] wl1[71] wl2[71] wl1[72] wl2[72] wl1[73] wl2[73] wl1[74] wl2[74] wl1[75] wl2[75] wl1[76] wl2[76] wl1[77] wl2[77] wl1[78] wl2[78] wl1[79] wl2[79] wl1[80] wl2[80] wl1[81] wl2[81] wl1[82] wl2[82] wl1[83] wl2[83] wl1[84] wl2[84] wl1[85] wl2[85] wl1[86] wl2[86] wl1[87] wl2[87] wl1[88] wl2[88] wl1[89] wl2[89] wl1[90] wl2[90] wl1[91] wl2[91] wl1[92] wl2[92] wl1[93] wl2[93] wl1[94] wl2[94] wl1[95] wl2[95] wl1[96] wl2[96] wl1[97] wl2[97] wl1[98] wl2[98] wl1[99] wl2[99] wl1[100] wl2[100] wl1[101] wl2[101] wl1[102] wl2[102] wl1[103] wl2[103] wl1[104] wl2[104] wl1[105] wl2[105] wl1[106] wl2[106] wl1[107] wl2[107] wl1[108] wl2[108] wl1[109] wl2[109] wl1[110] wl2[110] wl1[111] wl2[111] wl1[112] wl2[112] wl1[113] wl2[113] wl1[114] wl2[114] wl1[115] wl2[115] wl1[116] wl2[116] wl1[117] wl2[117] wl1[118] wl2[118] wl1[119] wl2[119] wl1[120] wl2[120] wl1[121] wl2[121] wl1[122] wl2[122] wl1[123] wl2[123] wl1[124] wl2[124] wl1[125] wl2[125] wl1[126] wl2[126] wl1[127] wl2[127] q1[0] q2[0] d1[0] d2[0] q1[1] q2[1] d1[1] d2[1] q1[2] q2[2] d1[2] d2[2] q1[3] q2[3] d1[3] d2[3] q1[4] q2[4] d1[4] d2[4] q1[5] q2[5] d1[5] d2[5] q1[6] q2[6] d1[6] d2[6] q1[7] q2[7] d1[7] d2[7] we1[0] clk1 we_en1 precharge1_n we2[0] clk2 we_en2 precharge2_n mux1[0] mux2[0] mux1[1] mux2[1] mux1[2] mux2[2] mux1[3] mux2[3] DP8TColumn_128R8B4M
.ends DP8TColumnBlock_128R8B4M1W

.subckt DP8TBlock_512x8_342A1WE clk1 clk2 a1[0] a2[0] a1[1] a2[1] a1[2] a2[2] a1[3] a2[3] a1[4] a2[4] a1[5] a2[5] a1[6] a2[6] a1[7] a2[7] a1[8] a2[8] vss vdd q1[0] q1[1] q1[2] q1[3] q1[4] q1[5] q1[6] q1[7] q2[0] q2[1] q2[2] q2[3] q2[4] q2[5] q2[6] q2[7] d1[0] d1[1] d1[2] d1[3] d1[4] d1[5] d1[6] d1[7] d2[0] d2[1] d2[2] d2[3] d2[4] d2[5] d2[6] d2[7] we1[0] we2[0]
Xrowperiph1 vss vdd clk1 a1[0] a1[1] a1[2] a1[3] a1[4] a1[5] a1[6] a1[7] a1[8] wl1[0] wl1[1] wl1[2] wl1[3] wl1[4] wl1[5] wl1[6] wl1[7] wl1[8] wl1[9] wl1[10] wl1[11] wl1[12] wl1[13] wl1[14] wl1[15] wl1[16] wl1[17] wl1[18] wl1[19] wl1[20] wl1[21] wl1[22] wl1[23] wl1[24] wl1[25] wl1[26] wl1[27] wl1[28] wl1[29] wl1[30] wl1[31] wl1[32] wl1[33] wl1[34] wl1[35] wl1[36] wl1[37] wl1[38] wl1[39] wl1[40] wl1[41] wl1[42] wl1[43] wl1[44] wl1[45] wl1[46] wl1[47] wl1[48] wl1[49] wl1[50] wl1[51] wl1[52] wl1[53] wl1[54] wl1[55] wl1[56] wl1[57] wl1[58] wl1[59] wl1[60] wl1[61] wl1[62] wl1[63] wl1[64] wl1[65] wl1[66] wl1[67] wl1[68] wl1[69] wl1[70] wl1[71] wl1[72] wl1[73] wl1[74] wl1[75] wl1[76] wl1[77] wl1[78] wl1[79] wl1[80] wl1[81] wl1[82] wl1[83] wl1[84] wl1[85] wl1[86] wl1[87] wl1[88] wl1[89] wl1[90] wl1[91] wl1[92] wl1[93] wl1[94] wl1[95] wl1[96] wl1[97] wl1[98] wl1[99] wl1[100] wl1[101] wl1[102] wl1[103] wl1[104] wl1[105] wl1[106] wl1[107] wl1[108] wl1[109] wl1[110] wl1[111] wl1[112] wl1[113] wl1[114] wl1[115] wl1[116] wl1[117] wl1[118] wl1[119] wl1[120] wl1[121] wl1[122] wl1[123] wl1[124] wl1[125] wl1[126] wl1[127] mux1[0] mux1[1] mux1[2] mux1[3] columnclk1 precharge1_n we_en1 DP8TRowPeriphery_3_4_2_wl1
Xrowperiph2 vss vdd clk2 a2[0] a2[1] a2[2] a2[3] a2[4] a2[5] a2[6] a2[7] a2[8] wl2[0] wl2[1] wl2[2] wl2[3] wl2[4] wl2[5] wl2[6] wl2[7] wl2[8] wl2[9] wl2[10] wl2[11] wl2[12] wl2[13] wl2[14] wl2[15] wl2[16] wl2[17] wl2[18] wl2[19] wl2[20] wl2[21] wl2[22] wl2[23] wl2[24] wl2[25] wl2[26] wl2[27] wl2[28] wl2[29] wl2[30] wl2[31] wl2[32] wl2[33] wl2[34] wl2[35] wl2[36] wl2[37] wl2[38] wl2[39] wl2[40] wl2[41] wl2[42] wl2[43] wl2[44] wl2[45] wl2[46] wl2[47] wl2[48] wl2[49] wl2[50] wl2[51] wl2[52] wl2[53] wl2[54] wl2[55] wl2[56] wl2[57] wl2[58] wl2[59] wl2[60] wl2[61] wl2[62] wl2[63] wl2[64] wl2[65] wl2[66] wl2[67] wl2[68] wl2[69] wl2[70] wl2[71] wl2[72] wl2[73] wl2[74] wl2[75] wl2[76] wl2[77] wl2[78] wl2[79] wl2[80] wl2[81] wl2[82] wl2[83] wl2[84] wl2[85] wl2[86] wl2[87] wl2[88] wl2[89] wl2[90] wl2[91] wl2[92] wl2[93] wl2[94] wl2[95] wl2[96] wl2[97] wl2[98] wl2[99] wl2[100] wl2[101] wl2[102] wl2[103] wl2[104] wl2[105] wl2[106] wl2[107] wl2[108] wl2[109] wl2[110] wl2[111] wl2[112] wl2[113] wl2[114] wl2[115] wl2[116] wl2[117] wl2[118] wl2[119] wl2[120] wl2[121] wl2[122] wl2[123] wl2[124] wl2[125] wl2[126] wl2[127] mux2[0] mux2[1] mux2[2] mux2[3] columnclk2 precharge2_n we_en2 DP8TRowPeriphery_3_4_2_wl2
Xcolumnblock vss vdd columnclk1 columnclk2 precharge1_n precharge2_n we_en1 we_en2 wl1[0] wl1[1] wl1[2] wl1[3] wl1[4] wl1[5] wl1[6] wl1[7] wl1[8] wl1[9] wl1[10] wl1[11] wl1[12] wl1[13] wl1[14] wl1[15] wl1[16] wl1[17] wl1[18] wl1[19] wl1[20] wl1[21] wl1[22] wl1[23] wl1[24] wl1[25] wl1[26] wl1[27] wl1[28] wl1[29] wl1[30] wl1[31] wl1[32] wl1[33] wl1[34] wl1[35] wl1[36] wl1[37] wl1[38] wl1[39] wl1[40] wl1[41] wl1[42] wl1[43] wl1[44] wl1[45] wl1[46] wl1[47] wl1[48] wl1[49] wl1[50] wl1[51] wl1[52] wl1[53] wl1[54] wl1[55] wl1[56] wl1[57] wl1[58] wl1[59] wl1[60] wl1[61] wl1[62] wl1[63] wl1[64] wl1[65] wl1[66] wl1[67] wl1[68] wl1[69] wl1[70] wl1[71] wl1[72] wl1[73] wl1[74] wl1[75] wl1[76] wl1[77] wl1[78] wl1[79] wl1[80] wl1[81] wl1[82] wl1[83] wl1[84] wl1[85] wl1[86] wl1[87] wl1[88] wl1[89] wl1[90] wl1[91] wl1[92] wl1[93] wl1[94] wl1[95] wl1[96] wl1[97] wl1[98] wl1[99] wl1[100] wl1[101] wl1[102] wl1[103] wl1[104] wl1[105] wl1[106] wl1[107] wl1[108] wl1[109] wl1[110] wl1[111] wl1[112] wl1[113] wl1[114] wl1[115] wl1[116] wl1[117] wl1[118] wl1[119] wl1[120] wl1[121] wl1[122] wl1[123] wl1[124] wl1[125] wl1[126] wl1[127] wl2[0] wl2[1] wl2[2] wl2[3] wl2[4] wl2[5] wl2[6] wl2[7] wl2[8] wl2[9] wl2[10] wl2[11] wl2[12] wl2[13] wl2[14] wl2[15] wl2[16] wl2[17] wl2[18] wl2[19] wl2[20] wl2[21] wl2[22] wl2[23] wl2[24] wl2[25] wl2[26] wl2[27] wl2[28] wl2[29] wl2[30] wl2[31] wl2[32] wl2[33] wl2[34] wl2[35] wl2[36] wl2[37] wl2[38] wl2[39] wl2[40] wl2[41] wl2[42] wl2[43] wl2[44] wl2[45] wl2[46] wl2[47] wl2[48] wl2[49] wl2[50] wl2[51] wl2[52] wl2[53] wl2[54] wl2[55] wl2[56] wl2[57] wl2[58] wl2[59] wl2[60] wl2[61] wl2[62] wl2[63] wl2[64] wl2[65] wl2[66] wl2[67] wl2[68] wl2[69] wl2[70] wl2[71] wl2[72] wl2[73] wl2[74] wl2[75] wl2[76] wl2[77] wl2[78] wl2[79] wl2[80] wl2[81] wl2[82] wl2[83] wl2[84] wl2[85] wl2[86] wl2[87] wl2[88] wl2[89] wl2[90] wl2[91] wl2[92] wl2[93] wl2[94] wl2[95] wl2[96] wl2[97] wl2[98] wl2[99] wl2[100] wl2[101] wl2[102] wl2[103] wl2[104] wl2[105] wl2[106] wl2[107] wl2[108] wl2[109] wl2[110] wl2[111] wl2[112] wl2[113] wl2[114] wl2[115] wl2[116] wl2[117] wl2[118] wl2[119] wl2[120] wl2[121] wl2[122] wl2[123] wl2[124] wl2[125] wl2[126] wl2[127] mux1[0] mux1[1] mux1[2] mux1[3] mux2[0] mux2[1] mux2[2] mux2[3] we1[0] we2[0] q1[0] q2[0] d1[0] d2[0] q1[1] q2[1] d1[1] d2[1] q1[2] q2[2] d1[2] d2[2] q1[3] q2[3] d1[3] d2[3] q1[4] q2[4] d1[4] d2[4] q1[5] q2[5] d1[5] d2[5] q1[6] q2[6] d1[6] d2[6] q1[7] q2[7] d1[7] d2[7] DP8TColumnBlock_128R8B4M1W
.ends DP8TBlock_512x8_342A1WE
Xtop clk1 clk2 a1[0] a2[0] a1[1] a2[1] a1[2] a2[2] a1[3] a2[3] a1[4] a2[4] a1[5] a2[5] a1[6] a2[6] a1[7] a2[7] a1[8] a2[8] vss vdd q1[0] q1[1] q1[2] q1[3] q1[4] q1[5] q1[6] q1[7] q2[0] q2[1] q2[2] q2[3] q2[4] q2[5] q2[6] q2[7] d1[0] d1[1] d1[2] d1[3] d1[4] d1[5] d1[6] d1[7] d2[0] d2[1] d2[2] d2[3] d2[4] d2[5] d2[6] d2[7] we1[0] we2[0] DP8TBlock_512x8_342A1WE
Vvss vss 0 0.0
Cq1[0] q1[0] 0 1e-14
Cq2[0] q2[0] 0 1e-14
Cq1[1] q1[1] 0 1e-14
Cq2[1] q2[1] 0 1e-14
Cq1[2] q1[2] 0 1e-14
Cq2[2] q2[2] 0 1e-14
Cq1[3] q1[3] 0 1e-14
Cq2[3] q2[3] 0 1e-14
Cq1[4] q1[4] 0 1e-14
Cq2[4] q2[4] 0 1e-14
Cq1[5] q1[5] 0 1e-14
Cq2[5] q2[5] 0 1e-14
Cq1[6] q1[6] 0 1e-14
Cq2[6] q2[6] 0 1e-14
Cq1[7] q1[7] 0 1e-14
Cq2[7] q2[7] 0 1e-14
Cq1[8] q1[8] 0 1e-14
Cq2[8] q2[8] 0 1e-14
Cq1[9] q1[9] 0 1e-14
Cq2[9] q2[9] 0 1e-14
Cq1[10] q1[10] 0 1e-14
Cq2[10] q2[10] 0 1e-14
Cq1[11] q1[11] 0 1e-14
Cq2[11] q2[11] 0 1e-14
Cq1[12] q1[12] 0 1e-14
Cq2[12] q2[12] 0 1e-14
Cq1[13] q1[13] 0 1e-14
Cq2[13] q2[13] 0 1e-14
Cq1[14] q1[14] 0 1e-14
Cq2[14] q2[14] 0 1e-14
Cq1[15] q1[15] 0 1e-14
Cq2[15] q2[15] 0 1e-14
Cq1[16] q1[16] 0 1e-14
Cq2[16] q2[16] 0 1e-14
Cq1[17] q1[17] 0 1e-14
Cq2[17] q2[17] 0 1e-14
Cq1[18] q1[18] 0 1e-14
Cq2[18] q2[18] 0 1e-14
Cq1[19] q1[19] 0 1e-14
Cq2[19] q2[19] 0 1e-14
Cq1[20] q1[20] 0 1e-14
Cq2[20] q2[20] 0 1e-14
Cq1[21] q1[21] 0 1e-14
Cq2[21] q2[21] 0 1e-14
Cq1[22] q1[22] 0 1e-14
Cq2[22] q2[22] 0 1e-14
Cq1[23] q1[23] 0 1e-14
Cq2[23] q2[23] 0 1e-14
Cq1[24] q1[24] 0 1e-14
Cq2[24] q2[24] 0 1e-14
Cq1[25] q1[25] 0 1e-14
Cq2[25] q2[25] 0 1e-14
Cq1[26] q1[26] 0 1e-14
Cq2[26] q2[26] 0 1e-14
Cq1[27] q1[27] 0 1e-14
Cq2[27] q2[27] 0 1e-14
Cq1[28] q1[28] 0 1e-14
Cq2[28] q2[28] 0 1e-14
Cq1[29] q1[29] 0 1e-14
Cq2[29] q2[29] 0 1e-14
Cq1[30] q1[30] 0 1e-14
Cq2[30] q2[30] 0 1e-14
Cq1[31] q1[31] 0 1e-14
Cq2[31] q2[31] 0 1e-14
Vvdd vdd_i 0 1.3
Rvdd vdd_i vdd 0.1
Vclk1 clk1_i 0 PWL(0.0s 0.0V 1e-08s 0.0V 1.02e-08s 1.3V 1.5000000000000002e-08s 1.3V 1.52e-08s 0.0V 2e-08s 0.0V 2.02e-08s 1.3V 2.5e-08s 1.3V 2.5199999999999997e-08s 0.0V)
Rclk1 clk1_i clk1 0.1
Vclk2 clk2_i 0 PWL(0.0s 0.0V 1e-08s 0.0V 1.02e-08s 1.3V 1.5000000000000002e-08s 1.3V 1.52e-08s 0.0V 2e-08s 0.0V 2.02e-08s 1.3V 2.5e-08s 1.3V 2.5199999999999997e-08s 0.0V)
Rclk2 clk2_i clk2 0.1
Va1[0] a1[0]_i 0 PWL(0.0s 0.0V 1.75e-08s 0.0V 1.77e-08s 1.3V)
Ra1[0] a1[0]_i a1[0] 0.1
Va1[1] a1[1]_i 0 PWL(0.0s 0.0V 1.75e-08s 0.0V 1.77e-08s 1.3V)
Ra1[1] a1[1]_i a1[1] 0.1
Va1[2] a1[2]_i 0 PWL(0.0s 0.0V 1.75e-08s 0.0V 1.77e-08s 1.3V)
Ra1[2] a1[2]_i a1[2] 0.1
Va1[3] a1[3]_i 0 PWL(0.0s 0.0V 1.75e-08s 0.0V 1.77e-08s 1.3V)
Ra1[3] a1[3]_i a1[3] 0.1
Va1[4] a1[4]_i 0 PWL(0.0s 0.0V 1.75e-08s 0.0V 1.77e-08s 1.3V)
Ra1[4] a1[4]_i a1[4] 0.1
Va1[5] a1[5]_i 0 PWL(0.0s 0.0V 1.75e-08s 0.0V 1.77e-08s 1.3V)
Ra1[5] a1[5]_i a1[5] 0.1
Va1[6] a1[6]_i 0 PWL(0.0s 0.0V 1.75e-08s 0.0V 1.77e-08s 1.3V)
Ra1[6] a1[6]_i a1[6] 0.1
Va1[7] a1[7]_i 0 PWL(0.0s 0.0V 1.75e-08s 0.0V 1.77e-08s 1.3V)
Ra1[7] a1[7]_i a1[7] 0.1
Va1[8] a1[8]_i 0 PWL(0.0s 0.0V 1.75e-08s 0.0V 1.77e-08s 1.3V)
Ra1[8] a1[8]_i a1[8] 0.1
Va2[0] a2[0]_i 0 PWL(0.0s 1.3V 1.75e-08s 1.3V 1.77e-08s 0.0V)
Ra2[0] a2[0]_i a2[0] 0.1
Va2[1] a2[1]_i 0 PWL(0.0s 1.3V 1.75e-08s 1.3V 1.77e-08s 0.0V)
Ra2[1] a2[1]_i a2[1] 0.1
Va2[2] a2[2]_i 0 PWL(0.0s 1.3V 1.75e-08s 1.3V 1.77e-08s 0.0V)
Ra2[2] a2[2]_i a2[2] 0.1
Va2[3] a2[3]_i 0 PWL(0.0s 1.3V 1.75e-08s 1.3V 1.77e-08s 0.0V)
Ra2[3] a2[3]_i a2[3] 0.1
Va2[4] a2[4]_i 0 PWL(0.0s 1.3V 1.75e-08s 1.3V 1.77e-08s 0.0V)
Ra2[4] a2[4]_i a2[4] 0.1
Va2[5] a2[5]_i 0 PWL(0.0s 1.3V 1.75e-08s 1.3V 1.77e-08s 0.0V)
Ra2[5] a2[5]_i a2[5] 0.1
Va2[6] a2[6]_i 0 PWL(0.0s 1.3V 1.75e-08s 1.3V 1.77e-08s 0.0V)
Ra2[6] a2[6]_i a2[6] 0.1
Va2[7] a2[7]_i 0 PWL(0.0s 1.3V 1.75e-08s 1.3V 1.77e-08s 0.0V)
Ra2[7] a2[7]_i a2[7] 0.1
Va2[8] a2[8]_i 0 PWL(0.0s 1.3V 1.75e-08s 1.3V 1.77e-08s 0.0V)
Ra2[8] a2[8]_i a2[8] 0.1
Vd1[0] d1[0]_i 0 1.3
Rd1[0] d1[0]_i d1[0] 0.1
Vd1[1] d1[1]_i 0 1.3
Rd1[1] d1[1]_i d1[1] 0.1
Vd1[2] d1[2]_i 0 1.3
Rd1[2] d1[2]_i d1[2] 0.1
Vd1[3] d1[3]_i 0 1.3
Rd1[3] d1[3]_i d1[3] 0.1
Vd1[4] d1[4]_i 0 1.3
Rd1[4] d1[4]_i d1[4] 0.1
Vd1[5] d1[5]_i 0 1.3
Rd1[5] d1[5]_i d1[5] 0.1
Vd1[6] d1[6]_i 0 1.3
Rd1[6] d1[6]_i d1[6] 0.1
Vd1[7] d1[7]_i 0 1.3
Rd1[7] d1[7]_i d1[7] 0.1
Vd1[8] d1[8]_i 0 1.3
Rd1[8] d1[8]_i d1[8] 0.1
Vd1[9] d1[9]_i 0 1.3
Rd1[9] d1[9]_i d1[9] 0.1
Vd1[10] d1[10]_i 0 1.3
Rd1[10] d1[10]_i d1[10] 0.1
Vd1[11] d1[11]_i 0 1.3
Rd1[11] d1[11]_i d1[11] 0.1
Vd1[12] d1[12]_i 0 1.3
Rd1[12] d1[12]_i d1[12] 0.1
Vd1[13] d1[13]_i 0 1.3
Rd1[13] d1[13]_i d1[13] 0.1
Vd1[14] d1[14]_i 0 1.3
Rd1[14] d1[14]_i d1[14] 0.1
Vd1[15] d1[15]_i 0 1.3
Rd1[15] d1[15]_i d1[15] 0.1
Vd1[16] d1[16]_i 0 1.3
Rd1[16] d1[16]_i d1[16] 0.1
Vd1[17] d1[17]_i 0 1.3
Rd1[17] d1[17]_i d1[17] 0.1
Vd1[18] d1[18]_i 0 1.3
Rd1[18] d1[18]_i d1[18] 0.1
Vd1[19] d1[19]_i 0 1.3
Rd1[19] d1[19]_i d1[19] 0.1
Vd1[20] d1[20]_i 0 1.3
Rd1[20] d1[20]_i d1[20] 0.1
Vd1[21] d1[21]_i 0 1.3
Rd1[21] d1[21]_i d1[21] 0.1
Vd1[22] d1[22]_i 0 1.3
Rd1[22] d1[22]_i d1[22] 0.1
Vd1[23] d1[23]_i 0 1.3
Rd1[23] d1[23]_i d1[23] 0.1
Vd1[24] d1[24]_i 0 1.3
Rd1[24] d1[24]_i d1[24] 0.1
Vd1[25] d1[25]_i 0 1.3
Rd1[25] d1[25]_i d1[25] 0.1
Vd1[26] d1[26]_i 0 1.3
Rd1[26] d1[26]_i d1[26] 0.1
Vd1[27] d1[27]_i 0 1.3
Rd1[27] d1[27]_i d1[27] 0.1
Vd1[28] d1[28]_i 0 1.3
Rd1[28] d1[28]_i d1[28] 0.1
Vd1[29] d1[29]_i 0 1.3
Rd1[29] d1[29]_i d1[29] 0.1
Vd1[30] d1[30]_i 0 1.3
Rd1[30] d1[30]_i d1[30] 0.1
Vd1[31] d1[31]_i 0 1.3
Rd1[31] d1[31]_i d1[31] 0.1
Vd2[0] d2[0]_i 0 0.0
Rd2[0] d2[0]_i d2[0] 0.1
Vd2[1] d2[1]_i 0 0.0
Rd2[1] d2[1]_i d2[1] 0.1
Vd2[2] d2[2]_i 0 0.0
Rd2[2] d2[2]_i d2[2] 0.1
Vd2[3] d2[3]_i 0 0.0
Rd2[3] d2[3]_i d2[3] 0.1
Vd2[4] d2[4]_i 0 0.0
Rd2[4] d2[4]_i d2[4] 0.1
Vd2[5] d2[5]_i 0 0.0
Rd2[5] d2[5]_i d2[5] 0.1
Vd2[6] d2[6]_i 0 0.0
Rd2[6] d2[6]_i d2[6] 0.1
Vd2[7] d2[7]_i 0 0.0
Rd2[7] d2[7]_i d2[7] 0.1
Vd2[8] d2[8]_i 0 0.0
Rd2[8] d2[8]_i d2[8] 0.1
Vd2[9] d2[9]_i 0 0.0
Rd2[9] d2[9]_i d2[9] 0.1
Vd2[10] d2[10]_i 0 0.0
Rd2[10] d2[10]_i d2[10] 0.1
Vd2[11] d2[11]_i 0 0.0
Rd2[11] d2[11]_i d2[11] 0.1
Vd2[12] d2[12]_i 0 0.0
Rd2[12] d2[12]_i d2[12] 0.1
Vd2[13] d2[13]_i 0 0.0
Rd2[13] d2[13]_i d2[13] 0.1
Vd2[14] d2[14]_i 0 0.0
Rd2[14] d2[14]_i d2[14] 0.1
Vd2[15] d2[15]_i 0 0.0
Rd2[15] d2[15]_i d2[15] 0.1
Vd2[16] d2[16]_i 0 0.0
Rd2[16] d2[16]_i d2[16] 0.1
Vd2[17] d2[17]_i 0 0.0
Rd2[17] d2[17]_i d2[17] 0.1
Vd2[18] d2[18]_i 0 0.0
Rd2[18] d2[18]_i d2[18] 0.1
Vd2[19] d2[19]_i 0 0.0
Rd2[19] d2[19]_i d2[19] 0.1
Vd2[20] d2[20]_i 0 0.0
Rd2[20] d2[20]_i d2[20] 0.1
Vd2[21] d2[21]_i 0 0.0
Rd2[21] d2[21]_i d2[21] 0.1
Vd2[22] d2[22]_i 0 0.0
Rd2[22] d2[22]_i d2[22] 0.1
Vd2[23] d2[23]_i 0 0.0
Rd2[23] d2[23]_i d2[23] 0.1
Vd2[24] d2[24]_i 0 0.0
Rd2[24] d2[24]_i d2[24] 0.1
Vd2[25] d2[25]_i 0 0.0
Rd2[25] d2[25]_i d2[25] 0.1
Vd2[26] d2[26]_i 0 0.0
Rd2[26] d2[26]_i d2[26] 0.1
Vd2[27] d2[27]_i 0 0.0
Rd2[27] d2[27]_i d2[27] 0.1
Vd2[28] d2[28]_i 0 0.0
Rd2[28] d2[28]_i d2[28] 0.1
Vd2[29] d2[29]_i 0 0.0
Rd2[29] d2[29]_i d2[29] 0.1
Vd2[30] d2[30]_i 0 0.0
Rd2[30] d2[30]_i d2[30] 0.1
Vd2[31] d2[31]_i 0 0.0
Rd2[31] d2[31]_i d2[31] 0.1
Vwe1[0] we1[0]_i 0 PWL(0.0s 1.3V 1.75e-08s 1.3V 1.77e-08s 0.0V)
Rwe1[0] we1[0]_i we1[0] 0.1
Vwe1[1] we1[1]_i 0 PWL(0.0s 1.3V 1.75e-08s 1.3V 1.77e-08s 0.0V)
Rwe1[1] we1[1]_i we1[1] 0.1
Vwe1[2] we1[2]_i 0 PWL(0.0s 1.3V 1.75e-08s 1.3V 1.77e-08s 0.0V)
Rwe1[2] we1[2]_i we1[2] 0.1
Vwe1[3] we1[3]_i 0 PWL(0.0s 1.3V 1.75e-08s 1.3V 1.77e-08s 0.0V)
Rwe1[3] we1[3]_i we1[3] 0.1
Vwe2[0] we2[0]_i 0 PWL(0.0s 1.3V 1.75e-08s 1.3V 1.77e-08s 0.0V)
Rwe2[0] we2[0]_i we2[0] 0.1
Vwe2[1] we2[1]_i 0 PWL(0.0s 1.3V 1.75e-08s 1.3V 1.77e-08s 0.0V)
Rwe2[1] we2[1]_i we2[1] 0.1
Vwe2[2] we2[2]_i 0 PWL(0.0s 1.3V 1.75e-08s 1.3V 1.77e-08s 0.0V)
Rwe2[2] we2[2]_i we2[2] 0.1
Vwe2[3] we2[3]_i 0 PWL(0.0s 1.3V 1.75e-08s 1.3V 1.77e-08s 0.0V)
Rwe2[3] we2[3]_i we2[3] 0.1

* Node initialization
.ic v(xtop.xrowperiph1.xcoldec.xaff[0]._dff_s)=0.0
.ic v(xtop.xrowperiph1.xcoldec.xaff[1]._dff_s)=0.0
.ic v(xtop.xrowperiph1.xrowdec.xpredec.xaff[0]._dff_s)=0.0
.ic v(xtop.xrowperiph1.xrowdec.xpredec.xaff[1]._dff_s)=0.0
.ic v(xtop.xrowperiph1.xrowdec.xpredec.xaff[2]._dff_s)=0.0
.ic v(xtop.xrowperiph1.xrowdec.xpredec.xaff[3]._dff_s)=0.0
.ic v(xtop.xrowperiph1.xrowdec.xpredec.xaff[4]._dff_s)=0.0
.ic v(xtop.xrowperiph1.xrowdec.xpredec.xaff[5]._dff_s)=0.0
.ic v(xtop.xrowperiph1.xrowdec.xpredec.xaff[6]._dff_s)=0.0
.ic v(xtop.xrowperiph2.xcoldec.xaff[0]._dff_s)=0.0
.ic v(xtop.xrowperiph2.xcoldec.xaff[1]._dff_s)=0.0
.ic v(xtop.xrowperiph2.xrowdec.xpredec.xaff[0]._dff_s)=0.0
.ic v(xtop.xrowperiph2.xrowdec.xpredec.xaff[1]._dff_s)=0.0
.ic v(xtop.xrowperiph2.xrowdec.xpredec.xaff[2]._dff_s)=0.0
.ic v(xtop.xrowperiph2.xrowdec.xpredec.xaff[3]._dff_s)=0.0
.ic v(xtop.xrowperiph2.xrowdec.xpredec.xaff[4]._dff_s)=0.0
.ic v(xtop.xrowperiph2.xrowdec.xpredec.xaff[5]._dff_s)=0.0
.ic v(xtop.xrowperiph2.xrowdec.xpredec.xaff[6]._dff_s)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[0])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[1])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[2])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[3])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[4])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[5])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[6])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[7])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[8])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[9])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[10])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[11])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[12])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[13])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[14])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[15])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[16])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[17])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[18])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[19])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[20])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[21])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[22])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[23])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[24])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[25])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[26])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[27])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[28])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[29])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[30])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1[31])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[0])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[1])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[2])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[3])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[4])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[5])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[6])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[7])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[8])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[9])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[10])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[11])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[12])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[13])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[14])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[15])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[16])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[17])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[18])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[19])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[20])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[21])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[22])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[23])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[24])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[25])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[26])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[27])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[28])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[29])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[30])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl1_n[31])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[0])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[1])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[2])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[3])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[4])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[5])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[6])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[7])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[8])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[9])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[10])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[11])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[12])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[13])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[14])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[15])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[16])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[17])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[18])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[19])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[20])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[21])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[22])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[23])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[24])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[25])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[26])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[27])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[28])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[29])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[30])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2[31])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[0])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[1])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[2])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[3])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[4])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[5])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[6])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[7])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[8])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[9])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[10])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[11])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[12])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[13])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[14])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[15])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[16])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[17])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[18])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[19])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[20])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[21])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[22])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[23])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[24])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[25])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[26])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[27])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[28])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[29])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[30])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].bl2_n[31])=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst0x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x0.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst0x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xarray.xinst1x0.xinst1x0.xinst1x0.xinst0x1.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.xinst0x1.xinst1x0.bit_n)=1.3
.ic v(xtop.xcolumnblock.xcolumn[0].xperiph1.xrw[0].xd_ff._dff_s)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xperiph1.xrw[1].xd_ff._dff_s)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xperiph1.xrw[2].xd_ff._dff_s)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xperiph1.xrw[3].xd_ff._dff_s)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xperiph1.xrw[4].xd_ff._dff_s)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xperiph1.xrw[5].xd_ff._dff_s)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xperiph1.xrw[6].xd_ff._dff_s)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xperiph1.xrw[7].xd_ff._dff_s)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xperiph1.xclkwe.xweff._dff_s)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xperiph2.xrw[0].xd_ff._dff_s)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xperiph2.xrw[1].xd_ff._dff_s)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xperiph2.xrw[2].xd_ff._dff_s)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xperiph2.xrw[3].xd_ff._dff_s)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xperiph2.xrw[4].xd_ff._dff_s)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xperiph2.xrw[5].xd_ff._dff_s)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xperiph2.xrw[6].xd_ff._dff_s)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xperiph2.xrw[7].xd_ff._dff_s)=0.0
.ic v(xtop.xcolumnblock.xcolumn[0].xperiph2.xclkwe.xweff._dff_s)=0.0
.save vss vdd
.save clk1 clk2
.save "a1[0]" "a1[1]" "a1[2]" "a1[3]" "a1[4]" "a1[5]" "a1[6]" "a1[7]" "a1[8]"
.save "d1[0]" "d1[1]" "d1[2]" "d1[3]" "d1[4]" "d1[5]" "d1[6]" "d1[7]"
.save "q1[0]" "q1[1]" "q1[2]" "q1[3]" "q1[4]" "q1[5]" "q1[6]" "q1[7]"
.save "we1[0]"
.save "a2[0]" "a2[1]" "a2[2]" "a2[3]" "a2[4]" "a2[5]" "a2[6]" "a2[7]" "a2[8]"
.save "d2[0]" "d2[1]" "d2[2]" "d2[3]" "d2[4]" "d2[5]" "d2[6]" "d2[7]"
.save "q2[0]" "q2[1]" "q2[2]" "q2[3]" "q2[4]" "q2[5]" "q2[6]" "q2[7]"
.save "we2[0]"
.save "xtop.mux1[0]" "xtop.mux1[1]"
.save "xtop.mux1[2]" "xtop.mux1[3]"
.save xtop.columnclk1 xtop.precharge1_n xtop.we_en1
.save "xtop.wl1[0]" "xtop.wl1[127]"
.save "xtop.mux2[0]" "xtop.mux2[1]"
.save "xtop.mux2[2]" "xtop.mux2[3]"
.save xtop.columnclk2 xtop.precharge2_n xtop.we_en2
.save "xtop.wl2[0]" "xtop.wl2[127]"
.save xtop.xrowperiph1.wl_en
.save "xtop.xrowperiph1.xrowdec.pd[0][0]"
.save "xtop.xrowperiph1.xrowdec.pd[0][1]"
.save "xtop.xrowperiph1.xrowdec.pd[0][2]"
.save "xtop.xrowperiph1.xrowdec.pd[0][3]"
.save "xtop.xrowperiph1.xrowdec.pd[0][4]"
.save "xtop.xrowperiph1.xrowdec.pd[0][5]"
.save "xtop.xrowperiph1.xrowdec.pd[0][6]"
.save "xtop.xrowperiph1.xrowdec.pd[0][7]"
.save "xtop.xrowperiph1.xrowdec.page[0]"
.save "xtop.xrowperiph1.xrowdec.page[1]"
.save "xtop.xrowperiph1.xrowdec.page[2]"
.save "xtop.xrowperiph1.xrowdec.page[3]"
.save "xtop.xrowperiph1.xrowdec.page[4]"
.save "xtop.xrowperiph1.xrowdec.page[5]"
.save "xtop.xrowperiph1.xrowdec.page[6]"
.save "xtop.xrowperiph1.xrowdec.page[7]"
.save "xtop.xrowperiph1.xrowdec.page[8]"
.save "xtop.xrowperiph1.xrowdec.page[9]"
.save "xtop.xrowperiph1.xrowdec.page[10]"
.save "xtop.xrowperiph1.xrowdec.page[11]"
.save "xtop.xrowperiph1.xrowdec.page[12]"
.save "xtop.xrowperiph1.xrowdec.page[13]"
.save "xtop.xrowperiph1.xrowdec.page[14]"
.save "xtop.xrowperiph1.xrowdec.page[15]"
.save xtop.xrowperiph2.wl_en
.save "xtop.xrowperiph2.xrowdec.pd[0][0]"
.save "xtop.xrowperiph2.xrowdec.pd[0][1]"
.save "xtop.xrowperiph2.xrowdec.pd[0][2]"
.save "xtop.xrowperiph2.xrowdec.pd[0][3]"
.save "xtop.xrowperiph2.xrowdec.pd[0][4]"
.save "xtop.xrowperiph2.xrowdec.pd[0][5]"
.save "xtop.xrowperiph2.xrowdec.pd[0][6]"
.save "xtop.xrowperiph2.xrowdec.pd[0][7]"
.save "xtop.xrowperiph2.xrowdec.page[0]"
.save "xtop.xrowperiph2.xrowdec.page[1]"
.save "xtop.xrowperiph2.xrowdec.page[2]"
.save "xtop.xrowperiph2.xrowdec.page[3]"
.save "xtop.xrowperiph2.xrowdec.page[4]"
.save "xtop.xrowperiph2.xrowdec.page[5]"
.save "xtop.xrowperiph2.xrowdec.page[6]"
.save "xtop.xrowperiph2.xrowdec.page[7]"
.save "xtop.xrowperiph2.xrowdec.page[8]"
.save "xtop.xrowperiph2.xrowdec.page[9]"
.save "xtop.xrowperiph2.xrowdec.page[10]"
.save "xtop.xrowperiph2.xrowdec.page[11]"
.save "xtop.xrowperiph2.xrowdec.page[12]"
.save "xtop.xrowperiph2.xrowdec.page[13]"
.save "xtop.xrowperiph2.xrowdec.page[14]"
.save "xtop.xrowperiph2.xrowdec.page[15]"
.save "xtop.xcolumnblock.xcolumn[0].bl1[0]" "xtop.xcolumnblock.xcolumn[0].bl1_n[0]"
.save "xtop.xcolumnblock.xcolumn[0].bl1[3]" "xtop.xcolumnblock.xcolumn[0].bl1_n[3]"
.save "xtop.xcolumnblock.xcolumn[0].bl2[0]" "xtop.xcolumnblock.xcolumn[0].bl2_n[0]"
.save "xtop.xcolumnblock.xcolumn[0].bl2[3]" "xtop.xcolumnblock.xcolumn[0].bl2_n[3]"
.save "xtop.xcolumnblock.xcolumn[0].xperiph1.muxbl[0]"
.save "xtop.xcolumnblock.xcolumn[0].xperiph1.muxbl_n[0]"
.save "xtop.xcolumnblock.xcolumn[0].xperiph1.xrw[0].bl_pd_g"
.save "xtop.xcolumnblock.xcolumn[0].xperiph1.xrw[0].bln_pd_g"
.save "xtop.xcolumnblock.xcolumn[0].xperiph2.muxbl[0]"
.save "xtop.xcolumnblock.xcolumn[0].xperiph2.muxbl_n[0]"
.save "xtop.xcolumnblock.xcolumn[0].xperiph2.xrw[0].bl_pd_g"
.save "xtop.xcolumnblock.xcolumn[0].xperiph2.xrw[0].bln_pd_g"
.save "xtop.xcolumnblock.xcolumn[0].bl1[28]" "xtop.xcolumnblock.xcolumn[3].bl1_n[28]"
.save "xtop.xcolumnblock.xcolumn[0].bl1[31]" "xtop.xcolumnblock.xcolumn[3].bl1_n[31]"
.save "xtop.xcolumnblock.xcolumn[0].bl2[28]" "xtop.xcolumnblock.xcolumn[3].bl2_n[28]"
.save "xtop.xcolumnblock.xcolumn[0].bl2[31]" "xtop.xcolumnblock.xcolumn[3].bl2_n[31]"
.save "xtop.xcolumnblock.xcolumn[0].xperiph1.muxbl[7]"
.save "xtop.xcolumnblock.xcolumn[0].xperiph1.muxbl_n[7]"
.save "xtop.xcolumnblock.xcolumn[0].xperiph1.xrw[7].bl_pd_g"
.save "xtop.xcolumnblock.xcolumn[0].xperiph1.xrw[7].bln_pd_g"
.save "xtop.xcolumnblock.xcolumn[0].xperiph2.muxbl[7]"
.save "xtop.xcolumnblock.xcolumn[0].xperiph2.muxbl_n[7]"
.save "xtop.xcolumnblock.xcolumn[0].xperiph2.xrw[7].bl_pd_g"
.save "xtop.xcolumnblock.xcolumn[0].xperiph2.xrw[7].bln_pd_g"
.options sparse method=gear
* take signal rise times as timestep
* take quarter of clock period as max time step
.tran 2e-10 3e-08 0.0 2.5e-09 uic
.end
